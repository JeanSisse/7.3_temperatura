library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_master is
	port(clk             : in  std_logic;
        address_a       : in  std_logic_vector(31 downto 2);
        enable_a        : in  std_logic;
        wbe_a           : in  std_logic_vector(3 downto 0);
        data_write_a    : in  std_logic_vector(31 downto 0);
        data_read_a     : out std_logic_vector(31 downto 0);

        address_b       : in  std_logic_vector(31 downto 2);
        enable_b        : in  std_logic;
        wbe_b           : in  std_logic_vector(3 downto 0);
        data_write_b    : in  std_logic_vector(31 downto 0);
        data_read_b     : out std_logic_vector(31 downto 0));
end; --entity ram     

architecture ram_master of ram_master is
signal enable_a_lo       : std_logic;
signal wbe_a_lo          : std_logic_vector(3 downto 0);
signal data_write_a_lo   : std_logic_vector(31 downto 0);
signal data_read_a_lo    : std_logic_vector(31 downto 0);
signal enable_b_lo       : std_logic;
signal wbe_b_lo          : std_logic_vector(3 downto 0);
signal data_read_b_lo    : std_logic_vector(31 downto 0);
signal enable_a_hi       : std_logic;
signal wbe_a_hi          : std_logic_vector(3 downto 0);
signal data_read_a_hi   : std_logic_vector(31 downto 0);
signal enable_b_hi       : std_logic;
signal wbe_b_hi          : std_logic_vector(3 downto 0);
signal data_read_b_hi    : std_logic_vector(31 downto 0);
signal address_a_reg     : std_logic_vector(31 downto 2);
signal address_b_reg     : std_logic_vector(31 downto 2);
signal enable_a_lo_256       : std_logic;
signal wbe_a_lo_256          : std_logic_vector(3 downto 0);
signal data_write_a_lo_256   : std_logic_vector(31 downto 0);
signal data_read_a_lo_256    : std_logic_vector(31 downto 0);
signal enable_b_lo_256       : std_logic;
signal wbe_b_lo_256          : std_logic_vector(3 downto 0);
signal data_read_b_lo_256    : std_logic_vector(31 downto 0);
signal enable_a_hi_256       : std_logic;
signal wbe_a_hi_256          : std_logic_vector(3 downto 0);
signal data_read_a_hi_256   : std_logic_vector(31 downto 0);
signal enable_b_hi_256       : std_logic;
signal wbe_b_hi_256          : std_logic_vector(3 downto 0);
signal data_read_b_hi_256    : std_logic_vector(31 downto 0);
begin
process(clk)
begin
if rising_edge(clk) then
	address_a_reg <= address_a;
	address_b_reg <= address_b;
	end if;
end process;
data_read_a <= data_read_a_lo when (address_a_reg < x"0001000"&"00") else
data_read_a_hi when ((address_a_reg >= x"0001000"&"00") and (address_a_reg < x"0002000"&"00")) else 
data_read_a_lo_256 when ((address_a_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_a_hi_256 when ((address_a_reg >= x"0003000"&"00") and (address_a_reg < x"0004000"&"00"));
data_read_b <= data_read_b_lo when (address_b_reg < x"0001000"&"00") else
data_read_b_hi when ((address_b_reg >= x"0001000"&"00") and (address_b_reg < x"0002000"&"00")) else
data_read_b_lo_256 when ((address_b_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_b_hi_256 when ((address_b_reg >= x"0003000"&"00") and (address_b_reg< x"0004000"&"00"));
enable_a_lo <= enable_a when (address_a < x"0001000"&"00") else '0';
enable_b_lo <= enable_b when (address_b < x"0001000"&"00") else '0';
enable_a_hi <= enable_a when ((address_a >= x"0001000"&"00") and (address_a < x"0002000"&"00")) else '0';
enable_b_hi <= enable_b when ((address_b >= x"0001000"&"00") and (address_b < x"0002000"&"00")) else '0';
enable_a_lo_256 <= enable_a when ((address_a >= x"0002000"&"00") and (address_a < x"0003000"&"00")) else '0';
enable_b_lo_256 <= enable_b when ((address_b >= x"0002000"&"00") and (address_b < x"0003000"&"00")) else '0';
enable_a_hi_256 <= enable_a when ((address_a >= x"0003000"&"00") and (address_a < x"0004000"&"00")) else '0';
enable_b_hi_256 <= enable_b when ((address_b >= x"0003000"&"00") and (address_b < x"0004000"&"00")) else '0';
wbe_a_lo <= wbe_a when  enable_a_lo='1' else x"0";
wbe_a_hi <= wbe_a when  enable_a_hi='1' else x"0";
wbe_b_lo <= wbe_b when  enable_b_lo='1' else x"0";
wbe_b_hi <= wbe_b when  enable_b_hi='1' else x"0";
wbe_a_lo_256 <= wbe_a when  enable_a_lo_256='1' else x"0";
wbe_a_hi_256 <= wbe_a when  enable_a_hi_256='1' else x"0";
wbe_b_lo_256 <= wbe_b when  enable_b_lo_256='1' else x"0";
wbe_b_hi_256 <= wbe_b when  enable_b_hi_256='1' else x"0";



ram_bit_0_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"88280C4C7B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"00160090920C04800904848262220277E05152B280780D407428E723C01E1400",
INIT_05 => X"0F001CC000890026105810941C5C06800E008057641E00473C40680D32330C00",
INIT_06 => X"82541A028D584E40CB0583CCA0100000161F84322000DA8C40F003C80030780E",
INIT_07 => X"BF70E1C3BBBB1138AF7F888025340C0888430047040FEE182CA00044BC5827C5",
INIT_08 => X"CAFC1F1F07F0FE1C94F65B11555EAFFC1C306758B24197ABCDA467F2C9CF9B32",
INIT_09 => X"4FFB4730000011420A61080800B6E0C464258094101606D5A47A2A2098B02000",
INIT_0A => X"446000304A0488111084048E082D0ED020119D35F900002FB00105C01036D800",
INIT_0B => X"1FA599581D3A9583C105A892112C04C0A898403120071501A6C32222068A3050",
INIT_0C => X"789E07A9E0789E07A9E0789E070CF0184F038850A21008E514845AB510D0106D",
INIT_0D => X"9A95E954868AD0E52273F4AC2180000808061C01C48B0F81380CE0F89E07A9E0",
INIT_0E => X"4001120055704FC4A1624487E2489024481224091282C4300942A19439481842",
INIT_0F => X"5D65C3E3F01F52FFC1E0013C1F801F52FFC1E0013C1F8090423D38A18E3B15C9",
INIT_10 => X"118796BE001F567FC1E0013C1F801F567FC1E0013C1F9085DFBF7E15C06101C5",
INIT_11 => X"7E30F00C0270F3751F1FD00FECBF7E25C0700463E17B2C7F811FD7ADECC381C0",
INIT_12 => X"4190626D6491063597F9177B956EF378D33E4030061341F077C571F8F885DFBF",
INIT_13 => X"7F328E3082636B2807FFD80FE00007E03F7207D3E03F9167184131B5C40FE647",
INIT_14 => X"EFA0CAE06101C53E3647D3F144FCDD22B81C0098E57D9081FCE8C8520C4DAE20",
INIT_15 => X"1ADF08DBF81846A540049707E0FE3307D3F141FFB45478040570EED41F4FE047",
INIT_16 => X"C189601208A1502B4AA5584B4068000019A80098120BCA4C617635C938574FF3",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"A800000000000000000902409024090240902409024090240902409024090240",
INIT_1A => X"08208208831042720EE38E38AAF9C4C704DAB63A6D58B3C10BAE8E789AA09424",
INIT_1B => X"7C3E1F0F87C3E1F0F82082082082082082082082082082082082082082082082",
INIT_1C => X"0003E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F8",
INIT_1D => X"0000000000000000000000000000000030F007FFFFFFFFFFFFFFFFFFFFFFF900",
INIT_1E => X"155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AEBDEBA0000000000000",
INIT_1F => X"7FD5545FF8000155087FC0155F7D168B55007BFDF45085168ABA002E82145085",
INIT_20 => X"55568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D7FFFE1000554214555",
INIT_21 => X"FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF7FFC00100800175555",
INIT_22 => X"0002E974BA5D5168A00A2D142155005142010FFAE820AAFF842AABAA2AE95545",
INIT_23 => X"AAFF803FFFF5D2A821550000000BA007FD55FF5D7FC0145007FD740055041541",
INIT_24 => X"FFF082EBDF455D5142000082E82145FFD17DFEFFFD168BFFF780000BA007FE8A",
INIT_25 => X"FE3F000000000000000000000000000000000000000000000AAFBEAA00007BFD",
INIT_26 => X"6F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEBDFD75D2AA8A80EA8E2",
INIT_27 => X"1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B68B551475FAF6D1C55",
INIT_28 => X"7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA0000542A0070071C50BAFEF",
INIT_29 => X"B8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A8010E004924874825D",
INIT_2A => X"EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0120155EA568E870BAE",
INIT_2B => X"7ABA497A82FFAFD2A82485FD2415A105C21451ED42A002545E055FFBE81D0BE8",
INIT_2C => X"00B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6A5C7E3DFFFE90B45B4",
INIT_2D => X"F45592E88A0AFE80A8B0A0000000000000000000000000000000000000000000",
INIT_2E => X"A1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE975EFAAAAB5E1AF3AABF",
INIT_2F => X"1CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB65F520EBE9EF67D7BE",
INIT_30 => X"034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EBC11472800752117082",
INIT_31 => X"968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F3142341D5DEEBEF55080",
INIT_32 => X"7D58AC448B69C30E02116220415A9540AA854140A0A2047F353AAF6C77F7F20D",
INIT_33 => X"56EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7C91565455C141E4188",
INIT_34 => X"F0000001FF0000001FF01EABC4B8014174FF7DA80F52FEDE6BE93172D7D625B5",
INIT_35 => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F",
INIT_36 => X"0000000000000000000000000000000000001FF0000001FF0000001FF0000001",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000100000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"CA1800080848B0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000010822C00803804000001999EF9C00040B0002000001000640200001018",
INIT_05 => X"08000000000100030008010468220A0004000000001000032000200002100800",
INIT_06 => X"8201961000060444010081002080000080820100000008004880000000284000",
INIT_07 => X"210C18306788C0089409800001140082000100010405000410A0000010082500",
INIT_08 => X"0A48903121780004C6000311555521F183060AC564BF818B5EDFDE0044600301",
INIT_09 => X"45B103200000140802234800000584000004808400020011A4581A2200002000",
INIT_0A => X"021000000800810400000402083000510000050020820036200005C00026C000",
INIT_0B => X"40000002000A008182200000002404400000000000010500008020A022220040",
INIT_0C => X"68064680646A0646A06468064690321503234204020018200404010784700404",
INIT_0D => X"C417C16004C0B838221090240180000801000C8800000190191064620646A064",
INIT_0E => X"6000000010200200802100022008100408020401020040100142200E0E08A20B",
INIT_0F => X"0021E300B000000781E00140018000000781E00140018000002430E30E0615C9",
INIT_10 => X"0000024E0000000781E00140018000000781E0014001908400005E11C0610000",
INIT_11 => X"3C30F00C000000155800D00000003E21C0700000000F00118000000468C381C0",
INIT_12 => X"40900004A400081401A0000004041218503E4030060000004804318008840000",
INIT_13 => X"01208C30800025200003D807E000000000725201600090461840001340002606",
INIT_14 => X"0F00C0E06100000012D2005100409520381C00000005920004C0C81200009A00",
INIT_15 => X"00120850B8180625400400000010711200510004B41478040000005548016000",
INIT_16 => X"40002002080000000804000A0000000011A000100208C008611430A000040250",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"0800000000000000000100401004010040100401004010040100401004010040",
INIT_1A => X"8A28A2AC8090C69606492492C09945235D5F7E2A5040B80E1C863A2958000500",
INIT_1B => X"DD6EB75BADD6EB75BAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A2",
INIT_1C => X"0002E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BA",
INIT_1D => X"00000000000000000000000000000000C0FFFFFFFFFFFFFFFFFFFFFFFFFFFC00",
INIT_1E => X"FE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5555550000000000000",
INIT_1F => X"D1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7AEBDF455D2EAABEFF7F",
INIT_20 => X"5000015500557DF45AAD1400BAA2AE801550051555EFF7AA95400552AAAABAFF",
INIT_21 => X"F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB5500517DF555D2EAAA105",
INIT_22 => X"5552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBAFFD540155557FD5400",
INIT_23 => X"10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAABAFF842ABEF5D517DF5",
INIT_24 => X"E105D2E954BAF7AE80010082A97410557FEABFFAAFBE8BEFAAD1575EF557FFFE",
INIT_25 => X"056A0000000000000000000000000000000000000000000005D7FFDF4500043F",
INIT_26 => X"BDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC51C7A2FBD5490BFD1C",
INIT_27 => X"4924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA974BAF7FFEFB45FFAA",
INIT_28 => X"DB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2080BEF495FC71D5412",
INIT_29 => X"FD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4002D082082AB8B6DBE",
INIT_2A => X"487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF78E021FF1471FDEAAF",
INIT_2B => X"FF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545A2DA3FB7DAAD4AAAAF",
INIT_2C => X"00547AB8F550A8010E00492487482FFFE82A85EBAE2FFC55554ADBD7A2FFC7BE",
INIT_2D => X"545AAFBF7400FBF9424F70000000000000000000000000000000000000000000",
INIT_2E => X"74AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E5400021EF005162BEF047FD5",
INIT_2F => X"225FF5843404547184164AA5D2EBEEB0A2D555410D3555714F8338AAAA1D0AE9",
INIT_30 => X"409000512AEABFFDF79DCBF755962010BDCBBC21455D7FEABEF75550ACBB7582",
INIT_31 => X"0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3FFEAAEB083BC1000FF8",
INIT_32 => X"BD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF801F8BA0C57740BDAA",
INIT_33 => X"DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF5D16BABAA3EBC3157A",
INIT_34 => X"0000000000000000000596EBEF55080034E0A592A4AD00FB863550229BCABEB7",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000100000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0812",
INIT_01 => X"A145A00810790848048044A54E404340404000720885800802000906E4910200",
INIT_02 => X"5C010802020408040C455850AA055254090541A111200A104A0000000908B510",
INIT_03 => X"182002200C00004485264A001214912803150020218808002440854288890550",
INIT_04 => X"210302048014100160806B08702010102722C9E0412200651102418214049492",
INIT_05 => X"88510910540008812C06010018204342A58A08011290A1120A81230240018DCA",
INIT_06 => X"47450000022480090000210002A54C282122040CC9082D530085224410AA4204",
INIT_07 => X"2101020423408900940C402A900011012D41D518044C10025000AA8A50043D00",
INIT_08 => X"214912534123010085008010141521F020409260000100A00004428808102010",
INIT_09 => X"519D12041551589141A539C42A4C9608080004801700D10100311820A848E0AA",
INIT_0A => X"0244C28C000002025A81AE3048321002A700200900160AE42CAA839AA90442C1",
INIT_0B => X"42300225604004D080251121D0000400880178044355940A498C400004A00545",
INIT_0C => X"4F240472404F240472404D240441200692022B41365E53340EC6940564D012D6",
INIT_0D => X"00000620500403080A919000038AD03001C5080D1108C1009001404524045240",
INIT_0E => X"02AA40AA902408000010002220040C000201030201200C818098402082020438",
INIT_0F => X"0080A0000140000002000140200A8000000200014020100280E469C698353000",
INIT_10 => X"000003400A800000020001402009400000020001402008700000000010000000",
INIT_11 => X"0004000000000081400004C00000000020000000008C000010A0000000100000",
INIT_12 => X"0000000680004188000400840080000000002000000000004810000001420000",
INIT_13 => X"0000000000003409280000000000000040025000030000000000001A05100000",
INIT_14 => X"000000000000000042900000A100000000000000008012A2000000000000D026",
INIT_15 => X"4420300000000000000000000010C010000098000000000000000105400002A0",
INIT_16 => X"126000808200505448342228120090554000E00000000000088000A000000000",
INIT_17 => X"004010040300C0300C0300C0100401004010040300C0300C0300C01004010240",
INIT_18 => X"0400004000040000C0200C0200C0200400004000040300C0300C0300C0100401",
INIT_19 => X"9FC0FC0FC1F81F81F800C0200C0200C0200400004000040000C0200C0200C020",
INIT_1A => X"0410411823A4301040B2CB2CBACB002009C6B860185AA1491B0E2863E8001100",
INIT_1B => X"4A25128944A25128941041041041041041041041041041041041041041041041",
INIT_1C => X"03F25128944A25128944A25128944A25128944A25128944A25128944A2512894",
INIT_1D => X"00000000000000000000000000000000F0F007FFFFFFFFFFFFFFFFFFFFFFFC07",
INIT_1E => X"415410AA8415555087BFFF55A2AA800BAFFAE9540008002AA000000000000000",
INIT_1F => X"FBEAABA5D7FE8B555551421455D0002145552EBFEBA007FC21EFA2FFD75EFAA8",
INIT_20 => X"2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F784155EFA2AEBDEAAA2",
INIT_21 => X"5D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BAA",
INIT_22 => X"55D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AAAAAAAAAAAFFD157410",
INIT_23 => X"FFA2D17DFEFF7800215500557DF55AA80001FFAA80001550055575EFFF840215",
INIT_24 => X"0AA082EAAB5500517DF555D042AA10A284154005D0015410085568A00FF80175",
INIT_25 => X"8A2A0000000000000000000000000000000000000000000005D00020AAAA8002",
INIT_26 => X"C51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA800AAFFAA9543A08003",
INIT_27 => X"0105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF49040017D5D20B8EAA007F",
INIT_28 => X"A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492AA8BC7EBDFEAFEFFD0",
INIT_29 => X"6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6FFEFB6D555578F7DB6",
INIT_2A => X"0155C51D0092A071555D5E3AE821D00001FF0871C016DBED1FDE90E3A497492B",
INIT_2B => X"8007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6DBE8F401D7B6A000147",
INIT_2C => X"00410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C5BE8555400550A3842",
INIT_2D => X"0AAF7AA954AA00042AAA20000000000000000000000000000000000000000000",
INIT_2E => X"21EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE975EF005560B55F7AA80",
INIT_2F => X"A8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BEABEF057D68F5F5A000",
INIT_30 => X"BFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D57DF55D7AABFF5428AC",
INIT_31 => X"D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002CA8AA80800020AAF7F",
INIT_32 => X"680800FFF7AAA155F595542455512A975455D3AA8A005500151FF0C57401E5F3",
INIT_33 => X"7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A2AA801455D7FE8BFFF",
INIT_34 => X"00000000000000000000C3BC1000FF8409000512AEABFF5D79FCAF774AE005BE",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000200000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380206",
INIT_01 => X"014C9A40408001683C0462C99E004B61404040028804A0080A000D16A0990A0C",
INIT_02 => X"4809A902031800444460589C66E331352180D468B8240E600C0081110B80ACD0",
INIT_03 => X"DA14C2210C0001D235834A0648D60528330006810A80881068A80C029CC56330",
INIT_04 => X"20886819A02740ECD2107364B37569100A04C1E01CA52010990240420E205A08",
INIT_05 => X"5831803532410000260E272058232259954369000A506912018CA582480038D1",
INIT_06 => X"8381A014000200AC2190ED0002ACD99881822144C5A409430682800046294140",
INIT_07 => X"218408142740E2C0948C3066500071913209CC8004640102D003999552083D20",
INIT_08 => X"00409231296AA180C2000110001521F0810A92E7402F00AB0016CA080C600111",
INIT_09 => X"41B112014D30E43802A76DD09905882B010605A01A4941010211088A2A43A399",
INIT_0A => X"4A12D9820880832264119D004860900104002008000F399606BC07998BA546AC",
INIT_0B => X"42522013604080D084A01001C8302D00008153000731C3000988C0040A224110",
INIT_0C => X"602406824068240602406224068920151203030032545B7404D7804566594796",
INIT_0D => X"080600E04C442068088590000999C8E84041086C001091009001406824060240",
INIT_0E => X"E6660599902600209021204A010E1C850C428521C208480021D842081A03E231",
INIT_0F => X"0090000003200000000010002008A00000000010002008038666928B28A65300",
INIT_10 => X"000801000A200000000010002009E0000000001000200A380000000000000000",
INIT_11 => X"0000000000000088000002D00000000000000000028010001620000000000000",
INIT_12 => X"0000008201021C88000048800280000000000000000004000010000003600000",
INIT_13 => X"8000000000041019980000000000000040802000068000000000020805B00000",
INIT_14 => X"0000000000000000C020000C8300000000000000008200AE000000000010402B",
INIT_15 => X"41003100000000000000000002008020000C3800000000000000012080001298",
INIT_16 => X"737420C20A01405468360022201185CCE0128410820000008088021C40A00008",
INIT_17 => X"2108721085218852188521885218852188521887210872108721087210872308",
INIT_18 => X"1086214872108621C852188421C852188421C852188721087210872108721087",
INIT_19 => X"26AA555AAB554AAB5561C852188421C852188421C85218842148721086214872",
INIT_1A => X"0410412881D0B0000092492480A981E063C638321450A08899A62C314A810508",
INIT_1B => X"EA753A9D4EA753A9D49249249249249249249249249249249249249241041041",
INIT_1C => X"BC4351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A9D4",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF82A",
INIT_1E => X"02AA00AA843DF55FFAA955EFA2D168B55557BEAA000055420000000000000000",
INIT_1F => X"5568A00087BE8BFFA2D155410AA8415555087BFFF55A2AA800BAFFAE95545080",
INIT_20 => X"D0002145552ABFEBA007FC21EF007FD75FFAA841541008002AB55AAAA955EF00",
INIT_21 => X"5D7FC0155005168B455D042AB45F7FFD741000042AA10AAAABFF5508003FF555",
INIT_22 => X"A5D7FC2010A2D1575FFF7AA975555D2E80145F78415545082EBDEAAA2FBEAABA",
INIT_23 => X"FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABFFF7FBEAB55F7AABDEB",
INIT_24 => X"B5555557DF55A2AEBDF555D2E954BA002EAAABA002A821EF5555554AA087BC01",
INIT_25 => X"203A000000000000000000000000000000000000000000000082E820BAA2FBEA",
INIT_26 => X"800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6FB7D5D7FEAA3808554",
INIT_27 => X"E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E1557D1475FAF45BEAA",
INIT_28 => X"AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2FBD55D7BE80004AA1E8",
INIT_29 => X"C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FFF5D0438140E2FA38B6",
INIT_2A => X"EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75D0A901FFFF801557D1",
INIT_2B => X"74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB455D20BDE00EBAAA8BC7",
INIT_2C => X"001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125FF002EADA921420871D",
INIT_2D => X"FFF5D7FEAABA0051400A20000000000000000000000000000000000000000000",
INIT_2E => X"75EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAAB55A28408145AAFFFF",
INIT_2F => X"D7145FBB8020A35D2ABEF55F7800015F087FEAA00007FEAB55FAD568AA2AFAE9",
INIT_30 => X"5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF55042AAAA007FD55558A7B",
INIT_31 => X"040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057968F575D003FF55F7D",
INIT_32 => X"52A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AAFFD5145FBAC9755F05",
INIT_33 => X"052ABFE10550415557085540000005156155FE90A8F5C082E974AAF7D57DF455",
INIT_34 => X"00000000000000000005500020AAF7FBFFFEF04552ABFFFF843FFE77C80825BC",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000100000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804002061080A284201081034809800A00230340007833522C82D04A16002",
INIT_01 => X"80439982183828490400050E12000340403008418984014902030106A0D10204",
INIT_02 => X"480108A000000000446418E01E80F00A41043118680402000800000009882390",
INIT_03 => X"0CA080210C0000408006480002001120260012603000000030808900888100F0",
INIT_04 => X"4403A609A055306B82C0705800CEE510082AC0A16B0350E3808041D03865D002",
INIT_05 => X"C0F20B36F0000901240626200820E26780E244A19A41E4020BAB06404001D312",
INIT_06 => X"434420151220118900806922406C3C7800201448DD9D2870020F228075A60715",
INIT_07 => X"2181000023480040840C001E180030032009700024641002C00187A440047C00",
INIT_08 => X"084830110160208004000001101121F220000260000100AA0004408000000001",
INIT_09 => X"519102063DF3E02B100B097407448F200A0209A041CA290102130C8800466478",
INIT_0A => X"8543D048006040064010E4007F62110105002002044007846124E0A00E0DC1EB",
INIT_0B => X"60020291404024808030512C40106D022203B1445810856A019400058F8404B5",
INIT_0C => X"052430D24305243052430D24304121A6921863013FD8807626EE000D64540284",
INIT_0D => X"28081080508104400A00800009B878680000880C1160410C90C143152430D243",
INIT_0E => X"81E0E18790012A00080102280800000202010102810020018098404110020004",
INIT_0F => X"0090000005E0200000001000200C6020000000100020000390E6C30830806204",
INIT_10 => X"000801000D20200000001000200EE0200000001000200A6A2000800000000000",
INIT_11 => X"8000000000000088000003B00100000000000000028000002EA0001000000000",
INIT_12 => X"80000082000251D80000C0044280000100000000000004000010000003282000",
INIT_13 => X"00002000000410121800040000000000408030000B8000100000020806F00000",
INIT_14 => X"0000100000000000C030000C9000008000000000008200FC000010000010403B",
INIT_15 => X"A500100000000100000000000200803000042E000200000000000120C0001590",
INIT_16 => X"30000800002400044934040AA231B63C20530801000410009889821040A00008",
INIT_17 => X"00401008000040300800004010000200C01000020040100802004030000002C0",
INIT_18 => X"000000C0300401008000000200C0100C01000020080000C030000000C0100802",
INIT_19 => X"325930C9A6CB261934C000200800004030040300800000020040100C03000000",
INIT_1A => X"8A28A2BD30264686668A28A2605145031C03F028000A1C2ED7831A2820244140",
INIT_1B => X"8D46A351A8D46A351AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A2",
INIT_1C => X"CFB068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D068351A",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF82B",
INIT_1E => X"54200000557FE10FFFBEAA10007FD7410FFAA97555082A800AA0000000000000",
INIT_1F => X"043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D168B55557BEAB45005",
INIT_20 => X"A8415555087BFFF55A2AA800BAFFAE9555508002AA000055574105D2A800AA00",
INIT_21 => X"087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAAA",
INIT_22 => X"0F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55A2AA955EF005568A00",
INIT_23 => X"AAA2FBD54BA080002145552ABFEAA007FC21EF007FD75FFAA8417410A2D14000",
INIT_24 => X"41000042AA10AAAABFF5508003FF55F7D568A00552EA8BEFA2AABDEAA087BEAA",
INIT_25 => X"50B800000000000000000000000000000000000000000000055042AB45F7FFD7",
INIT_26 => X"6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D5400F7A49057D08248",
INIT_27 => X"157428492E8008200043FE925571EFA380871C7028A28E3AF55F7A0925D7AADB",
INIT_28 => X"75C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA145",
INIT_29 => X"6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AAAEA8A9200249056D41",
INIT_2A => X"BE80004AAFEDB42028EBFBC2028BED152438AAA092492AAA4954281C0E2FB55B",
INIT_2B => X"FAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA007FC51C7007BD55D7",
INIT_2C => X"0041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEBAF7DF6AA00412EAABF",
INIT_2D => X"410FF84021EF0800154B20000000000000000000000000000000000000000000",
INIT_2E => X"AB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568A00FFFFEAA105D5155",
INIT_2F => X"955EF00042AAA25555410BA082E8201000043FE005D517DEBA0851574B2AAAEA",
INIT_30 => X"AAAA000804001FF005575408AA557FEB2FFAE975EF555168B55F7AA800BAF7AA",
INIT_31 => X"AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD568AA200557DE00AAA",
INIT_32 => X"07FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7D1550AAAA8002010F2",
INIT_33 => X"F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30800021EF55042AAAA0",
INIT_34 => X"000000000000000000008003FF55F7D5420BA5D2ABFEAAF7AEBDFF779A82AA43",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000200000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF0A0791B3FC1694378283C81FD996A091A32142007A336A20E03C040C002",
INIT_01 => X"A91FBDC4983088485C4A60000C24C26041280A00084000C8C212812EE2953231",
INIT_02 => X"C809AD5EB118E640A4F548FC011FF0002080000082ECC66609DB7DDDCB1FA036",
INIT_03 => X"4A120E4D3E4C90D294A31E824A52847A0B20640A88800000B8E0FD522885500E",
INIT_04 => X"001440849A2604001934800041110A71E2B068B110DB321C662AE22DC08A3448",
INIT_05 => X"370C14CA0E0800022446011C4E7F17907BEBD1AA65AE10571450DFC152522449",
INIT_06 => X"07319A109D129D450A846FE4E24C0305A1A5901C82416D05417118630839B88A",
INIT_07 => X"A5B56AD5A718C038AFFEA9FE39348C9204C389672407EE120EA5806E6C503AC5",
INIT_08 => X"C05896372728FF8C420619000003AFF4AD52A2C5D26F0EABCC96CD7AC4639902",
INIT_09 => X"5BD3571182080C000041080300F6F0C72221889C6FE20395A013282002B029F8",
INIT_0A => X"A23D203042444124098516CE0C2D13512410AD3CF8014005902DA6B2D1A4D810",
INIT_0B => X"645528937D5A85D3C4B0F883C10C24E0022B0E310612C2684CA16320A60A1185",
INIT_0C => X"288E3388E3208E3388E3288E330471904719C31438D04930ACE40FFD727C4304",
INIT_0D => X"8297A454544032252811E4AC2387F91008839C6CC413958D38C4E3208E3308E3",
INIT_0E => X"7FE0627FC25847C421516685844480204211200810028C38089AE00C894AA201",
INIT_0F => X"5D65E1E3C037E37FC3E0017C1F8037E37FC3E0017C1F900040261083080610CA",
INIT_10 => X"118796FE0037EA7FC3E0017C1F8037EA7FC3E0017C1F9300DFFFDE15D06101C5",
INIT_11 => X"BE34F00C0270F3754F1F8207FDBEBE25E0700463E17F3C7E054FF7BE6CD381C0",
INIT_12 => X"C090626DE40150459759573BBD6EF37D523E6030061341F07FC570F8FA00DFFF",
INIT_13 => X"6FE2AC3082636F301BFFFC07E00007E03F7263D383B7D1D6184131B7C1FEF64E",
INIT_14 => X"FFA0F0E06101C53E36E3D3EC84FDDDA8381C0098E57D923FDFC8D8120C4DBE0B",
INIT_15 => X"6FDF58DBF81C072540049707E0FE7323D3E43BFFF61478040570EED58F4F9397",
INIT_16 => X"00C108901822490448260224000040FC390250A2110B8ACC48B206A159A74FAB",
INIT_17 => X"08422080210882108C220842008821088230842208C20088210802308C2008C2",
INIT_18 => X"8422080230882108823080230842008C22084220842008C20080230802108C20",
INIT_19 => X"1092596D34924B2DA6884220842008821080230802108821084220842208C200",
INIT_1A => X"BEFBEFB7F7FE7EFEEE79E79EFAF2DDA73FBDCEDBFF9D3F0FDE0DB6DBF4208506",
INIT_1B => X"F77BBDDEEF77BBDDEEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"FED7BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF804",
INIT_1E => X"A800AAAAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF0000000000000",
INIT_1F => X"7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007FD7410FFAA97410082",
INIT_20 => X"A843DF55FFAA955EFA2D168B55557BEAB55005542000007FD74000055574BA5D",
INIT_21 => X"5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFFA",
INIT_22 => X"0F7D57FEBAFF80174BAAAD1555EF5555555550055574105D2A800AA00043FEBA",
INIT_23 => X"BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE95555080028A00A2FFFDE0",
INIT_24 => X"AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420BA5D2E821FFA2D5554",
INIT_25 => X"DFEF00000000000000000000000000000000000000000000000517FE10AAAAA8",
INIT_26 => X"D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC7010BEDF524AA5571F",
INIT_27 => X"1D74380851524BA5571D757DB6D5525EF555178F6D145178E00EBFBE8A101475",
INIT_28 => X"0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA147",
INIT_29 => X"92E8008200043FE925571EFA380871C7028B6AEBDF45B68A28B6DEBDF6DBEF1C",
INIT_2A => X"080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF55555057D1451524284",
INIT_2B => X"A552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45BEAA800AAFFAA9557D",
INIT_2C => X"0008517DE00AAAEA8A9200249056D4175C50920875FDA381C209256DFFDF420B",
INIT_2D => X"400F7FBC00BA55557DFF70000000000000000000000000000000000000000000",
INIT_2E => X"8A00AAFFEAA105D5155410FF84020AA0800154B2AAAA975FF5D7BC21EFF7FBD7",
INIT_2F => X"EABFF0051400A25551554BA0051400BA5551575EFF7D1401FF5D5568BE755556",
INIT_30 => X"AAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F78400145AAFFFFFEF5D7F",
INIT_31 => X"55421E75555400BA082E8201000043FE005D517DEBA0851574B2FFAABFF45FFA",
INIT_32 => X"7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF8002410FFD5575EF55",
INIT_33 => X"5D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7FFAE975EF555168B55F",
INIT_34 => X"000000000000000000000557DE00AAAAAAA000804001FF0055554088A557FEB2",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000C00000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000400322120040B313301C4389B2082",
INIT_01 => X"A74041CA38396849188160000C42424041000000090800090210090008110200",
INIT_02 => X"080108200C1000004465580000C0080100000000010432400800800009882050",
INIT_03 => X"080200010C234040842248600210812183806504488000103080014E88810000",
INIT_04 => X"0040504288A68210003120000000001002A0E8A910A072101000400A00203040",
INIT_05 => X"2800000400241801A52500094A02022014100128005004020010A1C044C02800",
INIT_06 => X"232000044084804914CA7C011AA3FC012122104CC0812D403280182308294000",
INIT_07 => X"2181020423488002940C0401D0480112000100004404004602447F8051223912",
INIT_08 => X"004812130160008304000000000021F020408264000108A00004400030400000",
INIT_09 => X"419102010104000A100348037F0584230A902A894008090343108802000FF407",
INIT_0A => X"B22D77C12052522400000400883011210000220006FC5FA400401484002447E0",
INIT_0B => X"60422291504420D084B0502044811428222300004611C57849A0150CA98A8561",
INIT_0C => X"1025B1025B0825B0825B1825B1112D8012D803003AD0413424E4014D627C0704",
INIT_0D => X"4404074040900B300A00810001A0021825E0886C0110916C96D15B0025B0025B",
INIT_0E => X"001E0800122100120499210A04A54652A12850962945180A14B44002CC020080",
INIT_0F => X"008ABA0030202100000001402068202100000001402067401026000000000031",
INIT_10 => X"00000341E8202800000001402068202800000001402062840000800000000000",
INIT_11 => X"8000000000000083D00052000100800000000000008CD0018400001200000000",
INIT_12 => X"800000069A48584000A0400000000005000000000000000048128D0002840000",
INIT_13 => X"80402000000034C1E000040000000000400FE000644000900000001A34000008",
INIT_14 => X"00003000000000004BA000112B0000880000000000807E80010010000000D1A4",
INIT_15 => X"0020250000040100000000000010CCE000198000020000000000010F80006028",
INIT_16 => X"0A728CA8C22540444924050CA9120603E0A2024048400010298432A002A00050",
INIT_17 => X"94E519465094A53946519425094A53946509425294E53946509425394E539625",
INIT_18 => X"425294E509425194E5294A519425094E5394A509465194A5294A519465094A52",
INIT_19 => X"3B1C618E38E38C31C71425294E53942519465294A53946509465394A50946519",
INIT_1A => X"8E38E39DB3B676F66EFBEFBEFAFBC5E73FC7F87A7D4ABFE7CFAFBE7BFA05004A",
INIT_1B => X"7F3F9FCFE7F3F9FCFE38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E3",
INIT_1C => X"6B23F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"00000000000000000000000000000000C0F007FFFFFFFFFFFFFFFFFFFFFFFC08",
INIT_1E => X"FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF0000000000000",
INIT_1F => X"AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFFBC0010AAD5574BA557",
INIT_20 => X"0557FE10FFFBEAA10007FD7410FFAA97400082A800AA08515555508043FE00F7",
INIT_21 => X"A2D5575EF55517FF55A2AA97400552AAAB45082E80155F7D1575EFFFAA955550",
INIT_22 => X"0FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD74000055574BA5D7FD7555",
INIT_23 => X"BAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000003DE1",
INIT_24 => X"B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE10AA803FE105D516AA",
INIT_25 => X"25FF000000000000000000000000000000000000000000000AAAEBDF45A28428",
INIT_26 => X"C7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49256DEB84104BAFFD15",
INIT_27 => X"B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE9756D145B401FFFFFF",
INIT_28 => X"DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A4904380824850381C5",
INIT_29 => X"851524BA5571D757DB6D5525EF555178F6DAAA495428412AAFB451C2A8017DE3",
INIT_2A => X"0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA2F1C50381471D74380",
INIT_2B => X"0A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D",
INIT_2C => X"00B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFFF1C7BD057D1C71FFE1",
INIT_2D => X"1FFAA84000AAFFD1401E70000000000000000000000000000000000000000000",
INIT_2E => X"75FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFDF55F78017400F78000",
INIT_2F => X"020AA0800154B2557FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2AAAA9",
INIT_30 => X"ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFFEAA105D5155410FF84",
INIT_31 => X"D5554B25551554BA0051400BA5551575EFF7D1401FF5D5568BE7AA80174AA082",
INIT_32 => X"AFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2AEA8A10082EA8BEFAA",
INIT_33 => X"557BC01EF55557DE00AA842AA0000516AABAFF8428BE7AAAEAAB55F78400145A",
INIT_34 => X"0000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000900000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0048201002842002C024500188000003000000003302300C018180006",
INIT_01 => X"020008402008404C042080000211024840000000080000080200010008110200",
INIT_02 => X"4801082248100000444008000080000041000000002222400800000009008010",
INIT_03 => X"0802010288A1484000020A400000002902006480088000003080040408810000",
INIT_04 => X"00004804890640004032030010000010008060E4100000140004500800403040",
INIT_05 => X"20000004004208016606010A0A20022000000000004000228010010080882000",
INIT_06 => X"030060004084004820906D311080020101000000008008011000000308290010",
INIT_07 => X"2100000023008002940C04000A4A010200018920646C10C50350002442003820",
INIT_08 => X"084812130160214204000000000121F000000244000100AA0004400920400000",
INIT_09 => X"419122810000081A00876882000590081100448A1000002350100CAA20002800",
INIT_0A => X"050280020100020400011640CC72602900044280028180242008069081244010",
INIT_0B => X"00200411508500B08805054C18024432A002400C99E410000080451100070014",
INIT_0C => X"05448054481544815448154481C22406A2406851201000200484950500F0145E",
INIT_0D => X"0144414A40000022880081511180036040044A013268E1205202480544805448",
INIT_0E => X"6000600010000020001102080102048102408120402800086098480008A20000",
INIT_0F => X"A2081210380021000001E003C0580021000001E003C042283426000000000021",
INIT_10 => X"00706801980028000001E003C0580028000001E003C044840000800009864038",
INIT_11 => X"80000330C00F0C0210807000010080000581C01C1C009201C000001200001607",
INIT_12 => X"8C2419101028D00020A2000000000005080082C180603A0E002A090404840000",
INIT_13 => X"8040204321188095F8000400061E001F800C202077C0009021908C4029F00008",
INIT_14 => X"00003009864038C10820201FAB000088026130071A00613E010011848322014F",
INIT_15 => X"6520350000640912058100F81C0108A0201FBA0002008239020F100880807BB8",
INIT_16 => X"114400C0002140144C2480200000040024A28400800044222980300CC4A0805C",
INIT_17 => X"2048120483204802008020082200812048120481200802008020081204812048",
INIT_18 => X"0880204812048020080200812048120080200802048320481204802008220080",
INIT_19 => X"2C208200010410400020C81200802008120C81204802008020C8120481200802",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000002A1050A",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"9840000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF818",
INIT_1E => X"5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04155550000000000000",
INIT_1F => X"AAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAAA97555F784174BAF7D",
INIT_20 => X"AAE955450055421FFFFFBC0010AAD5574BA557FFDFFF5555555EFAAFFFDFEFAA",
INIT_21 => X"A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00A",
INIT_22 => X"FA28000010552EBDE00007BEAAAAA2D14000008515555508043FE00F7AA97555",
INIT_23 => X"55557BD55FF00557FE10FFFBEAA10007FD7410FFAA97400082A800AAF7AE975F",
INIT_24 => X"B45082E80155F7D1575EFFFAA955555D51574AAAAFFD5545087FEAB455D516AB",
INIT_25 => X"7555000000000000000000000000000000000000000000000A2AA97400552AAA",
INIT_26 => X"9256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E1",
INIT_27 => X"B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7BFFF55FFA095482B6A4",
INIT_28 => X"2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF415",
INIT_29 => X"C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49003AFEFEBFBEAA001C",
INIT_2A => X"082485038F7A4905C7A28A070384120BDE100075EAA82BEDB470101C5B5057D1",
INIT_2B => X"5087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A101475D5400F7A490438",
INIT_2C => X"00AAA495428412AAFB451C2A8017DE3DF525FFFFA49756D495150492BEF1D255",
INIT_2D => X"A00555168A10002E9754D0000000000000000000000000000000000000000000",
INIT_2E => X"DF55F78017400F780001FFAA84000AAFFD1401E7FFAA97555A2AEA8A10AAD568",
INIT_2F => X"C00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215D557BF",
INIT_30 => X"028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7BC21EFF7FBD7400F7FB",
INIT_31 => X"FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2007FE8BFF080",
INIT_32 => X"D5155410FF84020AA0800154B2FF8402145A2AA954AA00043DE0000516AA10F7",
INIT_33 => X"005140000FFD140145007FE8BEF557BEAB55087FC215D555568A00AAFFEAA105",
INIT_34 => X"0000000000000000000AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"A140084000080048040100000202024040000000180800080200010048110204",
INIT_02 => X"080108020090000004655C000080000051000000002402400800000009008010",
INIT_03 => X"0002000100300C408422420002108108028065844880001030808D4288810000",
INIT_04 => X"0002584288A2C210003103001000001002A0E8C910A032541000090A00643040",
INIT_05 => X"2800080400645049A725010942220020140001A9005000004810A0C0044D2800",
INIT_06 => X"630400041404B141345A7C00426FFC01292214444081254102801A2308214004",
INIT_07 => X"21810204214080069408000008C3010200018920E06C0000021DFFA453263D32",
INIT_08 => X"084010110120018024000000000021F020408264000000080004400802400000",
INIT_09 => X"51B1004100040898128768820045142B0B902E895008080A1B13848A20002800",
INIT_0A => X"522920032052520400011641C460010D000000C8040100260008061081204010",
INIT_0B => X"4262229150012080102500211C81142880224000400411784920410C208514A4",
INIT_0C => X"0020000200002000020000200011000810008A55201000200484950004F0145E",
INIT_0D => X"40284301481509004885900101A0020964240109011890008011001020000200",
INIT_0E => X"0000200002210A320489000005A142D0A16850B6294D100A34B05242401340B4",
INIT_0F => X"00800008100001003C1FE00020080001003C1FE0002004401424008208041001",
INIT_10 => X"00000100080008003C1FE00020080008003C1FE000200080000001EA2F9EC000",
INIT_11 => X"01CB0FF3C000008000201000000081DA1F8FC0000080110080000002132C7E3F",
INIT_12 => X"3E6C00020040480040200000001004862CC19FCF81E000000010000200800000",
INIT_13 => X"004C11CF60001018000003F01FFE00004000000420800688E7B00008042000B8",
INIT_14 => X"000F251F9EC00000400004050002005D47E3F00000800084011607AD80004021",
INIT_15 => X"0000822406E5B85A3F830000000080000405000009AB87FB0000010000103000",
INIT_16 => X"1A768C68D260001448242704B912040002200640484000110104300042002018",
INIT_17 => X"B46D1B46D1B46D1B46D1B46D1B46D0B42D0B42D0B42D0B42D0B42D1B46D1B66D",
INIT_18 => X"46D1B42D0B42D0B42D0B42D1B46D1B46D1B46D1B42D0B42D0B42D0B42D0B42D0",
INIT_19 => X"200000000000000000346D1B46D1B46D0B42D0B42D0B42D0B46D1B46D1B46D1B",
INIT_1A => X"9E79E7B7F11E66C6FAD96D96520145052A1F5E2BD085122ED48F3AEB20840442",
INIT_1B => X"1F0F87C3E1F0F87C3E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"A6D4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF805",
INIT_1E => X"415555080000000087BEAA10F7803DE00FFAEBFFFF0800155FF0000000000000",
INIT_1F => X"80154105D7FC2145005155555F780155EFAAAEA8ABAAAFBFDE0055556AA005D0",
INIT_20 => X"87BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF552AA8AAA557FC0010F7",
INIT_21 => X"5D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF0",
INIT_22 => X"AAAAAA8B55F7D140010552E821EFAAAABDF555555555EFAAFFFDFEFAAAAAAB45",
INIT_23 => X"45557BE8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF5504000A",
INIT_24 => X"FFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F78402155AA8028A00A2D57FF",
INIT_25 => X"75D7000000000000000000000000000000000000000000000557BFDFFF55003D",
INIT_26 => X"FAE105D556AA10410E17555080E000280071E8A00EB8E3FE10F7AEBAFFF080A1",
INIT_27 => X"EA8AAA5571C2000FF8A17400557FC015514555757DFF8E175C7A2AAAAA82A2F1",
INIT_28 => X"FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF492",
INIT_29 => X"AF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A38492ABDE10EBDF7AF6DE3",
INIT_2A => X"5571FDFEF550E00082B6A0AFB55F7D1420104124821D7AAA0BDF6D415B575D7A",
INIT_2B => X"DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FFFFFFC7010BEDF524AA",
INIT_2C => X"00497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA001C2EA8A00F7800017",
INIT_2D => X"E00F7AEAABEF082E955450000000000000000000000000000000000000000000",
INIT_2E => X"7555A2AEA8A10AAD568A00555168A10002E9754D082E820BA08556AA00AAAABF",
INIT_2F => X"000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC21555D51575EFFFAA9",
INIT_30 => X"ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F78017400F780001FFAA84",
INIT_31 => X"843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215DA2FFE8ABA082",
INIT_32 => X"7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FFD540000000402145AA",
INIT_33 => X"5D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10AAAA975FF5D7BC21EFF",
INIT_34 => X"0000000000000000000007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000400000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000006",
INIT_01 => X"000009801830084C182060000C104268413C0A61590001D90213C10008110200",
INIT_02 => X"680108200010000054400C000080000041000000010002400800800009082011",
INIT_03 => X"0008000004002040000200100000000042800504488000103081880008C00000",
INIT_04 => X"00005042802A82100010030018000010000040C0100040140080040800003100",
INIT_05 => X"2000200400245001012100006002082000000000004000002010000040002000",
INIT_06 => X"2320400004040040144A7D000180020101000009808000000800001008210000",
INIT_07 => X"6100000021808000940800001800010200018B20206C01020200002441223C12",
INIT_08 => X"184010110120000004000000000061F000000244000081180004400000400000",
INIT_09 => X"4111002100040010008528820005100000900280000001000550860020002800",
INIT_0A => X"0080200520B23204000116404470900100402000000100242048025481024010",
INIT_0B => X"400000115040008002200000048034000002000000010712000000800F08A505",
INIT_0C => X"0000410004000041000400004100020000208201000000200404840284500016",
INIT_0D => X"00000120040000080000900201A0021924600088000000100100041000410004",
INIT_0E => X"60002000120002121C99024A00A14650A328519428651900142000000200A008",
INIT_0F => X"0000A20010200900000001400008200900000001400000001424008208041001",
INIT_10 => X"000002400820090000000140000820090000000140000A800000000000000000",
INIT_11 => X"0000000000000001500012000200800000000000000C10008400080200000000",
INIT_12 => X"0000000480004800002040000001000400000000000000004800010002800000",
INIT_13 => X"8041000000002401F80000000000000000025000274020800000001205D00808",
INIT_14 => X"004020000000000002900009AB00200800000000000012BA010100000000902E",
INIT_15 => X"652035000104000000000000001040100009BA000000000000000005400023B8",
INIT_16 => X"19028CA8D06540144C26832A1B0004000020024048400000090032A000000010",
INIT_17 => X"9425094250942509425094250942509425094250942509425094251946519465",
INIT_18 => X"4250942509425094250942519465194651946519465194651946519465194651",
INIT_19 => X"0800000000000000001465194651946519465194651946519425094250942509",
INIT_1A => X"34D34D1285B080201C92410480AB9A26667A46F345448020082E1C712A054008",
INIT_1B => X"1A0D068341A0D06834514514514514514514514514514514514514514D34D34D",
INIT_1C => X"2B60D069349A0D068341A4D268341A4D268341A0D069349A0D069349A0D06834",
INIT_1D => X"0000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF829",
INIT_1E => X"0155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA0000000000000",
INIT_1F => X"FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F7803DE00FFAEBFFFF080",
INIT_20 => X"780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555087BFDE00A2FBD7400F7",
INIT_21 => X"5D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA10F",
INIT_22 => X"A5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA557FC0010F78015410",
INIT_23 => X"45002EAAABA087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF780154A",
INIT_24 => X"E00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAABAF7D17FEBAA2AEBDF",
INIT_25 => X"8A92000000000000000000000000000000000000000000000AAFFE8A00552EBF",
INIT_26 => X"3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E",
INIT_27 => X"1FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E000280071E8A00EB8E",
INIT_28 => X"5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D556AA10410E17555087",
INIT_29 => X"571C2000FF8A17400557FC015514555757D5D71E8BEF147BFAE82A2DB555C71C",
INIT_2A => X"FFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A2AEADA38492EA8AAA5",
INIT_2B => X"2FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482B6A49256DEB84104BA",
INIT_2C => X"00A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D7000400155FFFBEDA8",
INIT_2D => X"B55FFAABDFEFF7D16AA000000000000000000000000000000000000000000000",
INIT_2E => X"20BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568BEF080402000F7AAA8",
INIT_2F => X"68A10002E9754D00517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00082E8",
INIT_30 => X"FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AEA8A10AAD568A005551",
INIT_31 => X"AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D51575EF555568BEF5D7",
INIT_32 => X"780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AAAE800AA552A97400A2",
INIT_33 => X"080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE00557BFDF55F78017400F",
INIT_34 => X"0000000000000000000A2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000800000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A14009821830284D182060000C10426840000000080000080200080000510204",
INIT_02 => X"0801080200100000046558040080000041000000002402400800000009008010",
INIT_03 => X"00020201040000D0842242024210810802006400088000003080054288C10000",
INIT_04 => X"0000400088020000003020002000001002A0E881108032100002000800203040",
INIT_05 => X"200000040000004924040108022000201000012800400010001081C040402000",
INIT_06 => X"030040040404804100006D2002A002012120004CC08125410200082308290000",
INIT_07 => X"2181020421408000940820001800010200018920206C01020200002440003C00",
INIT_08 => X"084010110120018004000000000021F020408264000000080004400800400000",
INIT_09 => X"511110010100008210010802004404230A000888400809000010042002002800",
INIT_0A => X"0000200000C04204000116404460910100082000040100240000000000004010",
INIT_0B => X"0AE22291404020902005002010000420A0200000400414684920410420200000",
INIT_0C => X"1120001200012001120011200011000090008840221000240484110000F05044",
INIT_0D => X"000803004C150100088480000980020000050001011890008011000120011200",
INIT_0E => X"000060001000020010010248040200010000800241000008009042404003E0BC",
INIT_0F => X"0080A00010202800000001402008202800000001402000000026008208041001",
INIT_10 => X"0000034008202100000001402008202100000001402002800000800000000000",
INIT_11 => X"8000000000000081400012000300000000000000008C10008400081000000000",
INIT_12 => X"8000000680001040002040000001000100000000000000004810000002800000",
INIT_13 => X"0001200000003408000004000000000040027000200020100000001A00000800",
INIT_14 => X"004010000000000042B00001000020800000000000801200000110000000D000",
INIT_15 => X"0000000001000100000000000010C030000100000200000000000105C0002000",
INIT_16 => X"03700080022100404D26A42EA01004002022000080000000018032A000A00010",
INIT_17 => X"0040100401004010040100401004010040100401004010040100400000000200",
INIT_18 => X"0000000000000000000000010040100401004010040100401004010040100401",
INIT_19 => X"0800000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"8A28A28D532A0CCC2A28A28A7AA344854A07F069CB8930AFD6A1AAA902A14148",
INIT_1B => X"6532994CA6532994CA28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A2",
INIT_1C => X"CC772B94CA6532994CA6572B95CAE532994CA6532995CAE572B94CA6532994CA",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF831",
INIT_1E => X"FEAABA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE100000000000000",
INIT_1F => X"8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA803DFFFAA843DF45FFF",
INIT_20 => X"80000000087BEAA10F7803DE00FFAEBFFFF0800155FF00042AB55FFD168B55AA",
INIT_21 => X"A2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE100",
INIT_22 => X"05555555EFF7FBC0145F78028A00A2D142155087BFDE00A2FBD7400F7FBFDFFF",
INIT_23 => X"FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555007FD741",
INIT_24 => X"EAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB55AAD168ABA002A975",
INIT_25 => X"8E00000000000000000000000000000000000000000000000557BE8BEF007FFD",
INIT_26 => X"38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E071D7AAFBEFB455D71F",
INIT_27 => X"42AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1E8B6D002090482B68E",
INIT_28 => X"D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D7000",
INIT_29 => X"2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD5410490A3DFD7F7A4821D7A2",
INIT_2A => X"410E175550071D54104951555D7EBF5C5155E3842AA00BED1421450871FFE00A",
INIT_2B => X"5BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82A2F1FAE105D556AA10",
INIT_2C => X"005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A38410E2ABD749516FB5",
INIT_2D => X"555A2FBFDF455D556AA000000000000000000000000000000000000000000000",
INIT_2E => X"8BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC01EFA2FFD7545AAAE97",
INIT_2F => X"AABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D56",
INIT_30 => X"EBFF45F78400155A2D57FE00552EA8A00082E820BA08556AA00AAAABFE00F7AE",
INIT_31 => X"D54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00FFFBD5400082",
INIT_32 => X"AD568A00555168A10002E9754D085155410085557555AAD557555A2802AA10FF",
INIT_33 => X"002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAFFAA97555A2AEA8A10A",
INIT_34 => X"0000000000000000000555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000008FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400986B830284D1820E0000C3642484000000008000008820009080A512220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"00080D4912E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"000048048002400048150300100002504230C8D9109032100020160880223000",
INIT_05 => X"220004440040080142020015001004A01200012840440000B01088C0005C2400",
INIT_06 => X"431018040014804920906C74B320020121210045408165445220082008211002",
INIT_07 => X"A5B1220421408004A56E840008B90D0200018B60A0650D450FC800644A0438A0",
INIT_08 => X"485816170760268E04000000000323F42C50826490640D28088445B0E0419003",
INIT_09 => X"41F1654100000818128728820024002B3B01AC9540080824CA13008820A02800",
INIT_0A => X"0000203600E06204000116C14474A3650048CE64E40100260048025481024810",
INIT_0B => X"08C32E915D9C208070042420180D24C8802000284007126A4D21262C20200404",
INIT_0C => X"31CA821CA831CA831CA821CA83165410E541085102000024040490A000D01056",
INIT_0D => X"812203360410110A4000840E3180021040465501011934A005101431CA821CA8",
INIT_0E => X"60006000101004A01811064B050204810240812241280D00200A08044290A088",
INIT_0F => X"482A01AAEC3602330CD2A02952DC3502330CB4A0318B41400024008208041011",
INIT_10 => X"0144C0155C3502330CD2A02952DC3602330CB4A0318B5600C587149B6D0141B0",
INIT_11 => X"083B6A51005956308D1E8202C436375908AA840AD4513437640F15245B455163",
INIT_12 => X"62F47B2872400044959BC42B1060F0D036B80B548523136C158878D8FE04E587",
INIT_13 => X"0A2699AAA3794392000D81852B0A050C224180062085134CD1719564E020C670",
INIT_14 => X"C50500D94C8121713C02B555101C90705D71009604140C0418CE0C378F0B2701",
INIT_15 => X"828E024D8C50965A40821568A06113801505010334AA73AA0666DAC20AD57400",
INIT_16 => X"123408C0822040544D248604B2100400100084008001D0113920060CDC06A27C",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"0080200802008020080200812048120481204812048120481204812048120481",
INIT_19 => X"0000000000000000002008020080200802008020080200802008020080200802",
INIT_1A => X"2082082815220A4A380000002A8313044020C0605885026853A1082100A00142",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000008208208",
INIT_1C => X"F070000000000000100800000000000000000004020000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF801",
INIT_1E => X"FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA0000000000000",
INIT_1F => X"2A801FFF7FFE8A10A28000000007FC2155F7D155545AA80001EFAAFBEAB45557",
INIT_20 => X"AFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2AEBFF45FFAEBFEAA00",
INIT_21 => X"FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEFA",
INIT_22 => X"5557FC2010002A80010A2842AAAA007BFFF4500042AB55FFD168B55AA8000010",
INIT_23 => X"EFFFD540000080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00557FF4",
INIT_24 => X"FEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021FF5D00154BAF7FBE8B",
INIT_25 => X"70AA000000000000000000000000000000000000000000000A2FFD741055003D",
INIT_26 => X"071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142ABDFC7F78E3FE28B6840",
INIT_27 => X"EBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007BC217DEBDB55555AA8E",
INIT_28 => X"AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92BEA",
INIT_29 => X"BDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA28A28BFF082ABAE10B6",
INIT_2A => X"080A175D708517DF7D497BC5028142A87000A28A2AA92007FF8F7D00042AB7DE",
INIT_2B => X"F5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00EB8E3FE10F7AEBAFFF",
INIT_2C => X"00B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E00B6DB6AA28A280001F",
INIT_2D => X"F55F7AABDEAAF784154BA0000000000000000000000000000000000000000000",
INIT_2E => X"01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBFFEF007BE8BFF5D2ABD",
INIT_2F => X"BDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BA087FC",
INIT_30 => X"AA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF080402000F7AAA8B55FFAA",
INIT_31 => X"7FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D5555FFAAA",
INIT_32 => X"AAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D2E95400A2AEA8A0000",
INIT_33 => X"FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA082E820BA08556AA00A",
INIT_34 => X"0000000000000000000FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000800000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702484000000008000008820009280A553231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"421A0A0012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"02004000890200001837830011998C31C09060DC104000102002140900003548",
INIT_05 => X"240000C400000001E404001F064000A00800000020480010A4100100001C2000",
INIT_06 => X"0300D800C1960C4400006E10B900020181840001008040057840001308212000",
INIT_07 => X"652428112180C03E8E5A2C800A3F018200418927E06686450FF8006460003A00",
INIT_08 => X"9840903525281D4F460409000000E3F08D1202C5C26A0719CC96CC7BF4629900",
INIT_09 => X"491175E10000041000C52882008600843001E09F0000002CF810200022302800",
INIT_0A => X"00002000030003040081164FC469227D2008CFE09A8180248009021091004810",
INIT_0B => X"00010C13499F01B33A00ACC0000F04F800000011800000000000433800000000",
INIT_0C => X"20CBC20CBC30CBC20CBC20CBC3065E1865E1000100000820040482B280504016",
INIT_0D => X"E7F3F01F40401C17E800C7FF3B80020000035780460124F16F06BC20CBC30CBC",
INIT_0E => X"00002200004005002001408400000000000000000000053A4096F80705FA0201",
INIT_0F => X"7B2C53F2FC16691DB587201EDDF4162B1DB527201EDDC46070241001000200F5",
INIT_10 => X"01D5CC9794162B1DB587201EDDF416691DB527201EDDD884272592D6246FC1B1",
INIT_11 => X"8E995D5A825DBA569F9FF02547068618CD3CC45B7863AE7EC00D4B122A67DF2A",
INIT_12 => X"CA5C33717461C045B5B182019473D19D7CCD856106F31A683621BDFC28800725",
INIT_13 => X"0A652CC8E3538BBA01624E51AA6C0469AC5493F5688532966471A9C5F6208C6C",
INIT_14 => X"41E1F5759001B4AA1853E6D5144AA9C914C8608D2724A4C4118D992B866E2FB1",
INIT_15 => X"825682D4A36C0B0B4B85112B2C4A05D3E6D5051893335EB0072AA85A4F9B7400",
INIT_16 => X"00800000082100544D248020000004001DC0800000010E7F70171401DE07EAD9",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0401004010040100401004000000000000000000000000000000000000000000",
INIT_19 => X"0800000000000000000040100401004010040100401004010040100401004010",
INIT_1A => X"249249120780800016A28A288028DCA30444409B054A88C5890486582A210108",
INIT_1B => X"32190C86432190C8641041041041041041041041041041041041041049249249",
INIT_1C => X"007592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2592C864",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF83E",
INIT_1E => X"0000AAAA843FE0008557DFFF0800020105D557FEAA00557DE100000000000000",
INIT_1F => X"AA8200000557DFFFF7AA80000082ABDF5508557DF45002ABDFFFF7803DE10AA8",
INIT_20 => X"07FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AAD5420000051555FFA2",
INIT_21 => X"F7FFE8A10A28000000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA0",
INIT_22 => X"05D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45FFAEBFEAA002A801FF",
INIT_23 => X"FFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA000028A1",
INIT_24 => X"BFF002ABDE00A2AABFE10082ABFFEF085542000000417555002A820AA08557DF",
INIT_25 => X"DE10000000000000000000000000000000000000000000000AAD155555A28428",
INIT_26 => X"BDFC7F78E3FE28B684070AABE803AE38145B78FD7000005010495B7AE921C517",
INIT_27 => X"547038145B505FFB6A487000005F7AFD7F7A482038002EBDF6D005B78F7D142A",
INIT_28 => X"2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00BED",
INIT_29 => X"BA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FFF1FDE821C003FE001C",
INIT_2A => X"F7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5D517DEAABEAEBFF7DE",
INIT_2B => X"5142082082005F7DFD7F7A482155BEF1E8B6D002090482B68E38FC7BE8A3DF7D",
INIT_2C => X"00B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FEF085F4703814001055",
INIT_2D => X"410007FEAA0055517DE000000000000000000000000000000000000000000000",
INIT_2E => X"FFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802AABA5D7FEAB45080015",
INIT_2F => X"FDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FEAB45F780020BA082EB",
INIT_30 => X"57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FFD7545AAAE97555A2FB",
INIT_31 => X"557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BAF7D1400BAFFD",
INIT_32 => X"7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA28428A105D7FEABEF55",
INIT_33 => X"087BD54AA550402145550000010087FFFF45F78402145F7D568BEF080402000F",
INIT_34 => X"0000000000000000000F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042604001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00020201926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"00104884880A4400403000004800027102A0E88110D83210642EA809C0203040",
INIT_05 => X"27000004004828032646000826080C201A008128044E00754010C9C192D82400",
INIT_06 => X"43000004080480492A946CE10320020121258044408125410270082308213800",
INIT_07 => X"A581424525408000AE2AA8002BC00D020003896020658FC4030000246E543AE5",
INIT_08 => X"4840101107200B80040210000002ABF02450A264002C80080004416800419000",
INIT_09 => X"4B531001000008001041080200B660E30B200C8840080A920651020002802800",
INIT_0A => X"0000203240E46204000516C04468C10100540034AC0100259001004010025010",
INIT_0B => X"04462E91440020905200A42209002420002800284002026A4D21758400000000",
INIT_0C => X"10000000000000010000000000000008000000000000002004040AA080504004",
INIT_0D => X"00000360401021280800E4000B800610C8410000A11210000000001000000000",
INIT_0E => X"6000600040D045E4195104D5854284A14250A12A512A8808289840084A020080",
INIT_0F => X"9E07A80948354B6E68982167061037496E683821670620681024000000000008",
INIT_10 => X"10B456587037496E689821670610354B6E6838216706220431961CA985D48094",
INIT_11 => X"186A91674011CE61403562274AA49CD594CF00039C7C414B6509DA22652138E5",
INIT_12 => X"3014780CC8604040424A5323845932E620295879818170304B2F5002C2043196",
INIT_13 => X"654B9104A328665603148895D44E0251142B42A3D8B2A5C8825194328A2E6A98",
INIT_14 => X"A6C6A465AA0091482382B17614F2202858EE300991415B45CD5306028F019451",
INIT_15 => X"08DC8047F17D1C7C3C02128E587D6A02B17605A130A4E8BF002258850AC5DC06",
INIT_16 => X"123508508220808048260604B2100C00022084809000D000393722A14000052E",
INIT_17 => X"284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A",
INIT_18 => X"84A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1",
INIT_19 => X"000000000000000000284A1284A1284A1284A1284A1284A1284A1284A1284A12",
INIT_1A => X"BAEBAEBFF6FEFEFEEEAAAAAAFBF7DDF77F9FBEFBFF9F3F0FDFCFBEFBF1228154",
INIT_1B => X"FD7EBF5FAFD7EBF5FAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAE",
INIT_1C => X"0077EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FA",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"57DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF0000000000000",
INIT_1F => X"7BEAB45552E80155AA802AB45AA843FE0008557DFFF0800020105D557FEAA005",
INIT_20 => X"82ABDF5508557DF45002ABDFFFF7803DE10AA80000AA087BD75EF087FFFFEF55",
INIT_21 => X"00557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAFFAE820AA5D55575550",
INIT_22 => X"FA2FBD7545FFD157555085140010F7AEAABFFAAD5420000051555FFA2AA82000",
INIT_23 => X"BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AAAEA8BF",
INIT_24 => X"EBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574BA557BE8A10A284154",
INIT_25 => X"ABD7000000000000000000000000000000000000000000000A2D155410F7FFFF",
INIT_26 => X"05010495B7AE921C517DE10A2DB50482147FFAF554971D0492E3F1C71C7BE8A2",
INIT_27 => X"1D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE803AE38145B78FD70000",
INIT_28 => X"A4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA1C7",
INIT_29 => X"45B505FFB6A487000005F7AFD7F7A482038AADF47092147FD257DFFD568A82FF",
INIT_2A => X"5D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000FFAAAFBFFBED5470381",
INIT_2B => X"24171EAA10B680124BAFFAAAFB45007BC217DEBDB55555AA8E071D7AAFBEFB45",
INIT_2C => X"00B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C20821C002AA92FFDF5748",
INIT_2D => X"010AAD157545F7AEA8B550000000000000000000000000000000000000000000",
INIT_2E => X"AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC00105D7BE8B55085142",
INIT_2F => X"BDEAAF784154BA5D5140145007BE8B55087BEAB555D04001EFF7AAA8B55F7802",
INIT_30 => X"FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007BE8BFF5D2ABDF55F7AA",
INIT_31 => X"AEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F780020BAA2FFD54105D7",
INIT_32 => X"AAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAAFBC0155085540000FF",
INIT_33 => X"5D042AA00F7FBD5410085568A10FF80020AAFFAABFF55087FC01EFA2FFD7545A",
INIT_34 => X"0000000000000000000F7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000CFFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"0002074F200904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000480488024000403000000000001002A0E881108032100002000800203040",
INIT_05 => X"200000040040080126060008020000201000012800400010001081C000402000",
INIT_06 => X"430000040004804920906C200220020121200044408125410200082308210000",
INIT_07 => X"A5A14285A15080008768A80008000D0200018B202067AF100A00002442043820",
INIT_08 => X"4850101105205380040000000000A7F42840A264920406080004400A00409002",
INIT_09 => X"411110010000080010010802000400230B000C88400808000211000002002800",
INIT_0A => X"0000203200E0620400011640446DA101004000002C0100240000000000004010",
INIT_0B => X"00422291400020900000002008002420002000004000026A4920410400000000",
INIT_0C => X"0000000000100000000000000100000000000000000000200404000000504004",
INIT_0D => X"0000022040100108080080000B80021040410000011010000000001000010000",
INIT_0E => X"0000600000000020181100400502048102408122412808082098400042020080",
INIT_0F => X"0040A100A42008000161C140000420080001C1C1400003201024000000000000",
INIT_10 => X"00022260042001000161C140000420010001C1C140001604E8084341CBA34048",
INIT_11 => X"2580E2B8802201014800C220A21829A302F1C024010C001124020C8C1A8A0396",
INIT_12 => X"0CA000048228404401004418012787124648157780120B8678C000801E04E808",
INIT_13 => X"072D04730000241000CB1325E78E0186030240000083B602398000120024ACA6",
INIT_14 => X"EF6F4163C480481506800004000CFD55196CB012481812049495C19400009001",
INIT_15 => X"800108B8FB61A0401200845594965000000400568D0CFB780055060500001001",
INIT_16 => X"123408408220000048240604B210040000008400800B0000090022A140068248",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"0481204812048120481204812048120481204812048120481204812048120481",
INIT_19 => X"0000000000000000002048120481204812048120481204812048120481204812",
INIT_1A => X"9E79E79FF3BEEEEEFE79E79EFAABCDA72E47F87BDF4EBAE7CFAFBEFB28200140",
INIT_1B => X"7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"FF83F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF83F",
INIT_1E => X"02ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA0000000000000",
INIT_1F => X"AE955455500155EF0804155EFAAD5554BA087FFFF55557BD54AAF7FBC01FFA28",
INIT_20 => X"A843FE0008557DFFF0800020105D557FEAA00557DE10A2AA801FFA28402000AA",
INIT_21 => X"552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400A",
INIT_22 => X"AA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF087FFFFEF557BEAB45",
INIT_23 => X"EF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA005568AB",
INIT_24 => X"555FFD168AAAFFAE820AA5D5557555002E80155A280000005D7FFDF4555517DF",
INIT_25 => X"0092000000000000000000000000000000000000000000000AAD1420AA087BD7",
INIT_26 => X"D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB4",
INIT_27 => X"E851FFB68402038AAAA955554900105FF0800175D7A2DB50482147FFAF554971",
INIT_28 => X"AAADB6D080A12410BE803AE38145B78FD7000005010495B7AE921C517DE10A2A",
INIT_29 => X"07FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2A0800BAE3F1C0092EB",
INIT_2A => X"B684070AA00516DABAA28402038B6803DE82F7F5D5410A2D568BC71C71D25D70",
INIT_2B => X"05D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D142ABDFC7F78E3FE28",
INIT_2C => X"00AADF47092147FD257DFFD568A82FFA4870BA555F5056D002A80155B6800001",
INIT_2D => X"145002AA8AAAAAFFC20000000000000000000000000000000000000000000000",
INIT_2E => X"00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFFF55FF84000AAAAFBC0",
INIT_2F => X"EAA0055517DE00A2AA955FFFF80020BAAAAA975450800001EF080417555A2FFC",
INIT_30 => X"0020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7FEAB45080015410007F",
INIT_31 => X"D56AB455D5140145007BE8B55087BEAB555D04001EFF7AAA8B555D557FE00A28",
INIT_32 => X"D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF803DE00FFD557400AA",
INIT_33 => X"082A80145F780020105D7BEAB45557BE8B45082EBFEBA082EBFFEF007BE8BFF5",
INIT_34 => X"0000000000000000000A2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000100000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"000440009282000001100000000000100220C8811080321000000228002A3000",
INIT_05 => X"200014C40000000100000000005C04A01000012A64400000145080C000422000",
INIT_06 => X"031042040804804100006EE4032002012120005540812540020008600831000A",
INIT_07 => X"21912244A14080008408880008000D0200018920206563000200002440003800",
INIT_08 => X"48501415032000800406180000002DF024408264000000080004400000430800",
INIT_09 => X"411100110000000010010802000400230A000880400808000450200000B02800",
INIT_0A => X"0000203000C042040001164044608101000000007C0100240000000000005810",
INIT_0B => X"0042229140002080000000200000040000200000400000684920000400000000",
INIT_0C => X"1000010000000000000000000100000800008000000000200404000010500004",
INIT_0D => X"00000260001001280000C4000300020000000000011010000000001000010000",
INIT_0E => X"400060000000000010010040040000000000000201000000000000004A000080",
INIT_0F => X"0000000000202100000000000000202100000000000004600024000000000008",
INIT_10 => X"0000000000202800000000000000202800000000000002000000800000000000",
INIT_11 => X"8000000000000000000002000100800000000000000000000400001200000000",
INIT_12 => X"80000000006000400080C0000000000D08120280000000000000000002000000",
INIT_13 => X"0040200000000010000004020010000000000000008000900000000000200008",
INIT_14 => X"0000308801400000000000040000008822110000000000040100100000000001",
INIT_15 => X"0000000004840717050000000000000000040000020000000000000000001000",
INIT_16 => X"023000000220000048240404A010040000008000000000000000020C40000008",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000200140",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"1420BAFF8000010082A954BA00003DFEF085155400F78428BEF0000000000000",
INIT_1F => X"843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD",
INIT_20 => X"AD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7AE95555A2FBE8BEFA2",
INIT_21 => X"5500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABAA",
INIT_22 => X"AA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FFA28402000AAAE95545",
INIT_23 => X"BA5D0015545AA843FE0008557DFFF0800020105D557FEAA00557DE10F7D1574A",
INIT_24 => X"0BAFFFFC20BAF7AEA8B45080417400FFFFC2145080015400AA802AA00AAAE800",
INIT_25 => X"DBFF00000000000000000000000000000000000000000000000516AA00A2AE80",
INIT_26 => X"50555412AA8ABAAADB40092E38E070280024904AA1C0438FD7005150438F78A2",
INIT_27 => X"A9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FFEDB55B6A080038E3DB",
INIT_28 => X"FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7E3A",
INIT_29 => X"68402038AAAA955554900105FF0800175D7E3FFEFBD70000124AA557FFDE10A2",
INIT_2A => X"1C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA38410038E38A2AE851FFB",
INIT_2B => X"0BE8E28A10AAA085082550A1057DBE803AE38145B78FD7000005010495B7AE92",
INIT_2C => X"001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A12410FFF1C017D14041040",
INIT_2D => X"B550855400AAF7AEBDFEF0000000000000000000000000000000000000000000",
INIT_2E => X"FF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA974AA0800020BA550028",
INIT_2F => X"57545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EFA2FBF",
INIT_30 => X"4020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7BE8B55085142010AAD1",
INIT_31 => X"002AAAAA2AA955FFFF80020BAAAAA975450800001EF080417555AAFFFDF45080",
INIT_32 => X"80015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7D17DF45007FE8AAA08",
INIT_33 => X"FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF7802AABA5D7FEAB450",
INIT_34 => X"00000000000000000005D557FE00A280020BAAAD140000A2AEBFFEF082A82010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000C00000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"0202115002BB10080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"2FE962000017102918900948514522CE09200C0D590569398ADBF8CC1E50E480",
INIT_05 => X"F05EA11E5600006B0800000038814B72A15B71D412E0AFD9C2990DA56FF0B55A",
INIT_06 => X"0640044150C025A0000000901A054F2C0A8030140BCC0460050690A95C8383D0",
INIT_07 => X"288500102F85203E8010D0AA9BC4800015001219D0550077373CAA8040006800",
INIT_08 => X"2064193920A2004B51400001414091EAA14881C0002701881B120203B7A80120",
INIT_09 => X"0409A02D965965200100104F2B00822512000000231520A024400800000ACCAA",
INIT_0A => X"0004B240028000342A00002FE00A3A1F06E649C005514AC40C082050010222D9",
INIT_0B => X"000A448C0082024AE50064B44000000000002A296AA000604838001980000000",
INIT_0C => X"044000440004400044000440004200022000200014808A02004200E540480212",
INIT_0D => X"0A80A5C8000102ED00440630004AD32400004000D58460018F6D3D8440004400",
INIT_0E => X"12AA28AA890BA00000024800480000000000000200802151025062C0BB400014",
INIT_0F => X"54E11C596A64003195933741477264003195555B418687E35836020814004049",
INIT_10 => X"99CF47DCB264003195933741597264003195555B4198843940076D296D0031F5",
INIT_11 => X"58486A556489347FE5F409CBC1362510695B6288743123C95251852041CD50A4",
INIT_12 => X"EAE2992046EB70026486035600CEC45CBCA809654B48163CCC895E1E043D4007",
INIT_13 => X"3A242DEA151848302BFD6D522B10C7EC71F6C1DB071D1216E078C4C1B1C74424",
INIT_14 => X"DAAABC982BE22267A2E2E4F44AA1DC5E37400C9EE1B7B638E8849D23C383298E",
INIT_15 => X"015998B28654565A003F0068E35352C1CAE48BFBF3A6C9B7B286B4DA8B93D037",
INIT_16 => X"009000040A8000452110A8442040D655602A102A0027E2C42320284086E6A2EE",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"1451451E96F2FC3C34F3CF3C2AC688AA263486D3260E34C0C3A7B451B0200000",
INIT_1B => X"7A7D1E9F47A7D1E9F4D14D14D14D14D14D14D14D14D14D14D14D14D145145145",
INIT_1C => X"0007D3E9F4FA7D3E8F47A3D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F4",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA0000000000000",
INIT_1F => X"80175EF0004000BA552A821FFFF8000010082A954BA00003DFEF085155400F78",
INIT_20 => X"2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D2E975EFF7D568BFFFF",
INIT_21 => X"AA8015400FF84001EF0000020AA5D00154005D043FF45555540000082EAABFFA",
INIT_22 => X"F5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555A2FBE8BEFA2843DE00",
INIT_23 => X"FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF557BEABE",
INIT_24 => X"4AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16ABFFFFAABFEAAFF84001",
INIT_25 => X"2092000000000000000000000000000000000000000000000FFFBE8BFF080017",
INIT_26 => X"38FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC",
INIT_27 => X"0925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E070280024904AA1C04",
INIT_28 => X"51420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB40092492",
INIT_29 => X"2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA410A1240055003FF6D55",
INIT_2A => X"BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC7557FC00BAE3AA9257DA",
INIT_2B => X"7F7AABAEAAF780051C70824851D7A2DB50482147FFAF554971D0492E3F1C71C7",
INIT_2C => X"00E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AABA08249756DF7D168BC",
INIT_2D => X"FFF552AAAAAA007BC00000000000000000000000000000000000000000000000",
INIT_2E => X"74AA0800020BA550028B550855400AAF7AEBDFEF08516AB55A2D16ABEFFFFBFD",
INIT_2F => X"A8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D04020AA002A955EFAAAA9",
INIT_30 => X"E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84000AAAAFBC0145002A",
INIT_31 => X"7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EF0800174BA002",
INIT_32 => X"85142010AAD157545F7AEA8B5500557DF45552A82000007BD74AAF7AEBDF455D",
INIT_33 => X"0804155FFF7D568B55FFAAAAABAFF8415545000015555A2FFC00105D7BE8B550",
INIT_34 => X"0000000000000000000AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000400000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"5295B6957FCBE0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"6DE90201BF90102103AF158E805428249851BFB2C106592088DBF8400A5055C2",
INIT_05 => X"403DA038338041EE341036BF36812841A19B68F40A807ED9C18114956FF081DB",
INIT_06 => X"00A0E2D7D3EAFF15800100FBFB333C1CBC303163670497AFF00291B3C0E20150",
INIT_07 => X"51C581123AEE54DE8008B719E61C10BBA5DAAFA9DDA1194D51E067BB00000000",
INIT_08 => X"0320A9392083056C2270E004400091181168C4D14002A110C902481FC0B42124",
INIT_09 => X"C51DFFC40C30E5F0182D0950190C0810BE00E9A76E4C6FFBE4700000B3038067",
INIT_0A => X"F7BC81C003C001674BB55B5FBB4BB4F26A19F70027CE86F047BEF19B6D94C1C1",
INIT_0B => X"0018CFC7429F326B9E822FFC00074D5A0AB033A3F330802966F74BFF8FCFB1F1",
INIT_0C => X"3EF3D3EF3D3EF3D3EF3D3EF3D3EF9E9F79E9E00185C44B91BC1740B7605040BE",
INIT_0D => X"CFEB69FF7A5F5AFFCCA787743FE67C21800367A28FC1AAF5CF6F3D3EF3D3EF3D",
INIT_0E => X"F99FD0678B87A0003000D8D02E00000000000000040025D3C21463D6BFF252D4",
INIT_0F => X"221ABD9CA854DFDD64A67D42C0F054DFDD64667D42C063E57A8F7B4594BB02C9",
INIT_10 => X"AA504801F054DFDD64A67D42C0F054DFDD64667D42C07237DFE5865F6D2BF232",
INIT_11 => X"8EAE7F5AB50D0806A9A2E0DFFF47DEDC496DA3181A0CC71440F9FBC3EFBB5AED",
INIT_12 => X"C3FC95949AEFF556EF9C75E7DCF1EB1B6E6FCDC87CB35FC94B36AECF3A33DFE5",
INIT_13 => X"AF5B6AAAE594A4C0DBFDAD94AA669809809FEFAF4157ADB55572CA527056E9C9",
INIT_14 => X"33F32ADD543430808BABAF50E1A5EB4BAEA45A250202FE0ADD39387F92B29382",
INIT_15 => X"523E865D4B1293AB6B90BF2F0E30EDEFAFD0B3FBD72E9E90D20A003FBEBF41AE",
INIT_16 => X"02F840000BCE0B6F67B3F845E017C833F6AAC02B002A2EFF22D4073DE83FB669",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9A69A6A4624C3434C0EBAEBA21B9001804F6E62029749701020B88A7CC0C0060",
INIT_1B => X"0D46A341A0D46A341A69AEBA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A6",
INIT_1C => X"00046A351A8D46A351A8D46A351A8D46A351A8D068341A0D068341A0D068341A",
INIT_1D => X"0000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA0000000000000",
INIT_1F => X"7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD17FFFF552EBFE00007",
INIT_20 => X"F8000010082A954BA00003DFEF085155400F78428BEFAAD168A000004020AA5D",
INIT_21 => X"0004000BA552A821FF5D00020BA552A82000552A821555D7FEAB55FF80175EFF",
INIT_22 => X"5AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EFF7D568BFFFF80175EF",
INIT_23 => X"55A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFFFFFDF4",
INIT_24 => X"4005D043FF45555540000082EAABFF00516AA10552E820BA007FEABEF0055555",
INIT_25 => X"AE920000000000000000000000000000000000000000000000000020AA5D0015",
INIT_26 => X"7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7",
INIT_27 => X"16AA381C0A07082497FEFB6D1451471EF007BD04920871F8FC7E3D56AB6DBEDB",
INIT_28 => X"7BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005150438F78A2DBFFBED",
INIT_29 => X"7D16ABFFE38E175EF1400000BA412E871FF550A00092492A850105D2A8015541",
INIT_2A => X"AADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5D7BFAEBA4920925EFF",
INIT_2B => X"2007FEDBD700515556DA2DF50492A2FFEDB55B6A080038E3DB50555412AA8ABA",
INIT_2C => X"000804050BA410A1240055003FF6D5551420101C2EAFBD7145B6AA2849248708",
INIT_2D => X"B550000175EFFFFBEAA000000000000000000000000000000000000000000000",
INIT_2E => X"AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFDFEFF7FBFFF55A2D16A",
INIT_2F => X"400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF5551555EF087FC200008516",
INIT_30 => X"A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800020BA550028B550855",
INIT_31 => X"7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002A955EF5D2E80010002",
INIT_32 => X"AFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FFD1575FF5504175EF5D",
INIT_33 => X"557FE8AAA000415410007BFFF450051555EFA2FBC0000A2FBFFF55FF84000AAA",
INIT_34 => X"00000000000000000000800174BA002E820105D003DFEF5D51420005D2ABFF45",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000CFFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"080BA868803F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"42016B0C401F58495C900A4859552A611D9A640F5903B2388004004C08A06008",
INIT_05 => X"7008000E0E508C01C28640000801133060E0032801E0202000991B708280B501",
INIT_06 => X"560000000022229A60B048048120FF040000000002C44D620F0228454C838100",
INIT_07 => X"58800A001D4033A004904087F9E3901218050018024110D6771C1F90C2856828",
INIT_08 => X"3020A82929A807B3731021400058C020000A9729400D10100420480202AC2140",
INIT_09 => X"0419002D86184A01018030430700802541420440022030041A814A0080064C1F",
INIT_0A => X"0000F0CA8428642430080438408A510185A200000045C18C0E0000A0820500B9",
INIT_0B => X"311324AA2373088479105D044A1022000001835C0C30C2E21480349D00100202",
INIT_0C => X"000C2000C2000C2000C2000C2000610006100100180A8062026000DC425C0301",
INIT_0D => X"10108003C00021002046088B5001FB3650D89844703657083080C2800C2000C2",
INIT_0E => X"007E281F840C00284A17210001060D8306C18360C1380A0260CB980840080810",
INIT_0F => X"9BBEF8E50B041029075982BF3873041029079982BF39748AA0AC800014804032",
INIT_10 => X"79BFD7F7F3041029075982BF3E73041029079982BF3F632C5F96D3C11555D5D7",
INIT_11 => X"A595405FC7F1CFEBC7586C4100A53162B47FD7E39FFEECE1598702345156AEA4",
INIT_12 => X"FE037ACFB88083A99E06271BB0CA207DFDD5920057E0B001B0EBCC79932C5F96",
INIT_13 => X"2A002DD51B6F7FC4A411D1E8D44517F14EAFE36E55150016EA8DB73E39464006",
INIT_14 => X"C30351452A13D55CFFA76E928E3891F148B30399F5FB7F28C800DFA06F5DF5CA",
INIT_15 => X"57DFEAEF1005475F1D1F608819CF0EE76E12C824ADD9089715F25FAF9DB84953",
INIT_16 => X"34041A41A0000010180C02801680460FC900052FA10DC0006DA4881C110155AC",
INIT_17 => X"60D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8",
INIT_18 => X"0D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D83",
INIT_19 => X"00000000000000000020D8360D8360D8360D8360D8360D8360D8360D8360D836",
INIT_1A => X"8A28A2891182C8A82E0820825945DF675C0770B9E11807E54587BEF8B0000000",
INIT_1B => X"2552A954AA5128944AAAA28A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A2",
INIT_1C => X"000128944A25128944A25128944A25128944A25128944A25128944A25128944A",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E954000000000000000",
INIT_1F => X"D568B55080028B55002E82000087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD",
INIT_20 => X"87FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA087FFFFFFFFFBFDF45AA",
INIT_21 => X"0051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE000",
INIT_22 => X"00804154BA55042ABEF5D7FD75FFAAD540145AAD168A000004020AA5D7BE8B45",
INIT_23 => X"10557FD7545FF8000010082A954BA00003DFEF085155400F78428BEFAA800000",
INIT_24 => X"000552A821555D7FEAB55FF80175EF5D00020105D2A97400082E95555085168A",
INIT_25 => X"24280000000000000000000000000000000000000000000005D00020BA552A82",
INIT_26 => X"E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A9",
INIT_27 => X"FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147FFFFFFFFFBFDFC7EBF5",
INIT_28 => X"003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092087",
INIT_29 => X"C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AADF6DB7DE3F5FAFC708",
INIT_2A => X"F78A2DBFFA28407038140410492550A2ABC7497BD25FFAADF4516DBED16AA381",
INIT_2B => X"8002E9557D1C516FA28417BD5545E38E070280024904AA1C0438FD7005150438",
INIT_2C => X"00550A00092492A850105D2A80155417BEFB6DEB8E175FF5D0E0500049209742",
INIT_2D => X"FEF552E974AA082A820AA0000000000000000000000000000000000000000000",
INIT_2E => X"DFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFFFFFFFFFFDFEFF7FBFF",
INIT_2F => X"AAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AA557FF",
INIT_30 => X"FFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D16ABEFFFFBFDFFF552A",
INIT_31 => X"FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087FC2000FFD56AB45A2F",
INIT_32 => X"50028B550855400AAF7AEBDFEFA280154BA550400000552AA8B45087FC01EFA2",
INIT_33 => X"5D2E974000804154BA082A975EF5D517DEAA007BD5545AAAA974AA0800020BA5",
INIT_34 => X"00000000000000000005D2E80010002A954005D2A82155087FFFFEFAAAA975EF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000400000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000010228001000000000000000000024001620280000000000354200004008",
INIT_04 => X"00016200001310090090004840004152C7208802590000388000004C08006000",
INIT_05 => X"7008000E0200000000000000000100302000000000E02000009900000000B100",
INIT_06 => X"00000000000000100000000000001B040000000002C42010010200004C838100",
INIT_07 => X"E0050A040041593104004500480090080A011202201400204204018000000000",
INIT_08 => X"30E409080188000021A0000100004082A140102B4020109801A4CE0037100100",
INIT_09 => X"00000005861840000000004301000B000000000001C1C0000000000000020C01",
INIT_0A => X"0000B0C0000000101400040C0408100000000000004540800000000000000099",
INIT_0B => X"000010000800011000000000000000000000BC0007C00008092C800080000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"08000EC0000000000000000010004B2000000000000000000000000000000000",
INIT_0E => X"0006280180040000000000000000000000000000000000000000000000000001",
INIT_0F => X"4451B81A70AB3006BA0011400760AB3006BA0011400680F02096834820000000",
INIT_10 => X"04082248A0AB3006BA0011400160AB3006BA0011400084C780687DBA82800808",
INIT_11 => X"796E80A00802301BC0A7531EDD98E73B02800804620D030F873EB49F30B80112",
INIT_12 => X"0000002044F091A860700FF9198AA115D5DA37F7A80C8A3604001C0664C78068",
INIT_13 => X"51AC9000000000314E01F9F30198600631448410A2A8D64800000081B0A936B0",
INIT_14 => X"0303842281C80A23004411AD661891F15148A4420804241526D6000000000985",
INIT_15 => X"35F3D282000C6C5456C84850F61050C411AD6284FDA861682805A04A1046B2E0",
INIT_16 => X"00000000000000000000000000004600C0013800003088004202304366A4A9D3",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"86186186851046260A9A69A6039045DD1F863808633005010063A20C90000000",
INIT_1B => X"930984C26130984C261861861869A61861861861869A61861861861861861861",
INIT_1C => X"0000984C26130984C26130984C26130984C26130984C26130984C26130984D26",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BA0000000000000",
INIT_1F => X"FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082",
INIT_20 => X"87FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7FFFFFFFFFFFFFFFFF7",
INIT_21 => X"080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA0",
INIT_22 => X"FF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFFFFFBFDF45AAD568B55",
INIT_23 => X"00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AAF7FFFFFF",
INIT_24 => X"B55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB55A2FFFDFEF5D2EBFE",
INIT_25 => X"04AA000000000000000000000000000000000000000000000AAFFFDF45A2D16A",
INIT_26 => X"FDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA00001",
INIT_27 => X"FFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7FFFFFFFFFFFFFFFF7FB",
INIT_28 => X"00001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92EBF",
INIT_29 => X"3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7F1F8FD7AAD16AB4500",
INIT_2A => X"087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D000000010087FFDFC7E",
INIT_2B => X"DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6DBEDB7FFEF552AB8E38",
INIT_2C => X"00B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E284971F8FC7AAD56DB6",
INIT_2D => X"FEF552E954AA0004000AA0000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFFFFFFFFFFFFFFFFFFFD",
INIT_2F => X"175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00557FF",
INIT_30 => X"56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FBFFF55A2D16AB550000",
INIT_31 => X"0402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AAF7FBFDFEFF7D",
INIT_32 => X"FFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7FFFFFFF552AA8BEF08",
INIT_33 => X"08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA0008516AB55A2D16ABEFF",
INIT_34 => X"0000000000000000000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000800000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"0001E6000053300B00D0005800000000000000407B0004BB830004DC3D01E000",
INIT_05 => X"F0FF433EFE022001C81080001101F977E0201C409BE1F10623BB000A100CF300",
INIT_06 => X"0F00100002E22EB440012C809B2FFF7C8E8840155FDC0000010E40087D8787A1",
INIT_07 => X"3B800000000000000008407FC800B0000000100600040000C205FF91C000F800",
INIT_08 => X"28C0B0300020852000002101554021F000000000000000090492260200002000",
INIT_09 => X"00000007BEFBC010002008FF7F00000000010018A81000041C401000004FFDFF",
INIT_0A => X"0002B7C0000008000000200000200A0C004408C2007D5FC800000240001227FB",
INIT_0B => X"000000000000000000000000800800A400000000000000008000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000800080000000",
INIT_0D => X"001000000100000020000800101FFB6000000000000000000000000000000000",
INIT_0E => X"07FE29FF800C00000001002040000000000000020480002E42429C0000080000",
INIT_0F => X"4D4E180010040000400000001E60040000400000001E6010003C000000000030",
INIT_10 => X"000094B1E0040000400000001E60040000400000001E60804000000400000000",
INIT_11 => X"02000000000033628000100100000004000000006170C0008001000004000000",
INIT_12 => X"000000295810000000A100020614148002000000000004307CC3CC0000804000",
INIT_13 => X"2000000000014AC000120200000000003F0D800020100000000000A4B0020000",
INIT_14 => X"0C0C00000000002E2D000001006204040000000005786C004000000000052580",
INIT_15 => X"0A0C0939BEE1810080200000E0CE0EC000010020000000000000AE8A00002002",
INIT_16 => X"8040400400C08080000000000049F6FFC0100000000000008008008000400010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000200",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C30C320624C1090D0F3CF3CD038001801C10000804482A60D09008269020010",
INIT_1B => X"86432190C86432190CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C3",
INIT_1C => X"000432190C86432190C86432190C86432190C86432190C86432190C86432190C",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"4174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804020100000000000000",
INIT_1F => X"FFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA000",
INIT_20 => X"87FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFFFFF",
INIT_21 => X"552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA0",
INIT_22 => X"FFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFFFFFFFFFFFF7FBFDFFF",
INIT_23 => X"EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA007FFFFF",
INIT_24 => X"FEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDFEFF7D56AB450000021",
INIT_25 => X"5000000000000000000000000000000000000000000000000F7FFFFFFFFFFFFD",
INIT_26 => X"FFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA08000",
INIT_27 => X"FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428087",
INIT_29 => X"FFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFFFFFFFEFF7FBFFFFF55",
INIT_2A => X"B6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AABEDF6FABAEBFFFFFFFF",
INIT_2B => X"7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7EBF5E8B550000071EF",
INIT_2C => X"00FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AAA497FFFFFFF7FBF8FC",
INIT_2D => X"FFF5D2A954AA0800174100000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410A2FFF",
INIT_30 => X"BFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFFFDFEFF7FBFFFEF552E",
INIT_31 => X"FFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00AAFFFFFFFFFF",
INIT_32 => X"2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAAD16AB450804174AAFF",
INIT_33 => X"087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA557FFDFEFF7FBFFF55A",
INIT_34 => X"0000000000000000000F7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"1094EC681244819000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"0001E6000053300F01D4587800446194F49020107F0012BBC00202DC3823EA82",
INIT_05 => X"F0F807BFFE000120080002341881F3FFF012412A9FE1E01013BF09404050F300",
INIT_06 => X"08808210996035A000006EC2E04FFFFC0A0000101FFE4036450E08247F878703",
INIT_07 => X"003400812A156C002822987FC830F40134CC74D002016612DE87FFE004008040",
INIT_08 => X"02348D2D00080C0C53400044114000000D022640B42406808790055043A82824",
INIT_09 => X"080AC707FEFBC110008420F7FF388B70A20389346FE8000580200800008FDFFF",
INIT_0A => X"4636FFC00080013029811240444A82422A828C03BC7D7FC15025B1AB6E85A7FF",
INIT_0B => X"2019480E63180855A492712CC01C49C20201BFE45FF0C004041DA2218A8A3151",
INIT_0C => X"648A3648A3648A3648A3648A366451B2451B210018C241102068006C620C0388",
INIT_0D => X"80050094104431200090080C621FFBE0008A94641165448C80C103648A3648A3",
INIT_0E => X"9FFEADFF8050250010030165290008800440022201082401A002000C48000201",
INIT_0F => X"48A004A6C0D2820302C005A83480D1820302A009B02B101390C0CB2830816202",
INIT_10 => X"8904831400D1820302C005A83480D2820302A009B02B021A85C0941150013180",
INIT_11 => X"8834600024D052C1051E0B92D400360520202682C19024B6164E300448510140",
INIT_12 => X"4093E22A2012418A9D1D44ADD9E0F174103820101C0B8160D5516259FA1A85C0",
INIT_13 => X"8AA288209E615100280DA0052000C5006402000206C55144104D510CC1B0D640",
INIT_14 => X"D50020C04023033C52009144231D902818100C90058010361AC808126C88660D",
INIT_15 => X"2386454988140600C0181500A13E830011008B0374007000B4E0CD00024500A0",
INIT_16 => X"0224004002000000703804008001F7FFF01B982B01258088C008CC41198A1220",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"0000000000000000002008020080200802008020080200802008020080200802",
INIT_1A => X"BEFBEFBFF7FEFEFFFE79E79FFFF7CFF77FBFFEFBFF9F7E0FDF9EFEFBF0000000",
INIT_1B => X"FF7FBFDFEFF7FBFDFEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000100000000000000",
INIT_1F => X"FFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080",
INIT_20 => X"7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAF",
INIT_22 => X"FFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFFFFFFFFFFFFFFFFFFEF",
INIT_23 => X"AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFF",
INIT_24 => X"FFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFFFFFFFBFDFEF5D2A954",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA00000",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAF7F",
INIT_29 => X"FFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFFFFFFFFFFFFFFDFEF55",
INIT_2A => X"082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA002A95400087FFFFFFF",
INIT_2B => X"FF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA",
INIT_2C => X"00E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50BA557FFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0000020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAFFFFF",
INIT_30 => X"FFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E",
INIT_31 => X"2E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410087FFFFFFFFF",
INIT_32 => X"7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7FBFFFFF552E954BA00",
INIT_33 => X"5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA557FFFFFFFFFFFDFEFF",
INIT_34 => X"0000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"8632CA211E4491D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"24B000808800040439245B221373581F97B0A8D1040F92000F42000047A00E58",
INIT_05 => X"0107C4410008816B105036B4180C000811E9BF2844021B1004045E4249500449",
INIT_06 => X"0111C2D50A46AE45281502E4A2200081ADA0E054402365774611E047020008E0",
INIT_07 => X"80BD5AA4BF5C91F840C1710010344DB9A808FDFF3DE0313014A2007540401804",
INIT_08 => X"EA212D6D481ADF0CE47CA21544009007A64EBD64049D028B93D9561A48F60276",
INIT_09 => X"0E48D500400015805060040080A2A0F4A82381B4000A0905A0283800AA500200",
INIT_0A => X"4E700838460402635019FBFE7FCA13520F8AAD050402204090090319A5002004",
INIT_0B => X"040F4A944B1AA313C0022AA0011C0DC0002800134000000849BCC3240A8A7151",
INIT_0C => X"70AA070AA070AA070AA070AA072550385503800500001840000C80B410014088",
INIT_0D => X"0A9CA0D458D131652A154CAC6B600085080B14004D1594832824A070AA070AA0",
INIT_0E => X"C00044000A1EC1C44140D101A54280A14050A028500A84F02842A24C594A0687",
INIT_0F => X"59E0C4E6C256690581800F1C3E82562B0581200F1C3F08145602280402080448",
INIT_10 => X"AB8581B602562B0581800F1C3E8256690581200F1C3F1238473F121000613383",
INIT_11 => X"0E1050083750B3E4275F829547008600C030374361FA2CEE046D48122C438100",
INIT_12 => X"C012A66F61154C019511628756231018500C00203E138061565160782238473F",
INIT_13 => X"AA612C0096C37B00D1724801A0009C606D1221D104553096004B61BCC1128C4C",
INIT_14 => X"41E0F0600035842E7601C2C4AC68A98810080AA825A890225189980254CDE608",
INIT_15 => X"637E00D0A1080301401C390320188321C2C0B13890105800D520AF94870B012A",
INIT_16 => X"22F110111B281A54753AA004002601001918008C10912A4440B24E8B58234A89",
INIT_17 => X"0882208822088220882208822088220882208822088220882208822088220882",
INIT_18 => X"8020080200802008020080200802008020080200802208822088220882208822",
INIT_19 => X"8000000001FFFFFFFFC802008020080200802008020080200802008020080200",
INIT_1A => X"9E79E7BFF3FEFEBEEEFBEFBEFBEFDFEF7F47F8FBEF5EB7E6CFEFBEFBE8289144",
INIT_1B => X"7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"0003F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000000000000000000",
INIT_1F => X"FFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFF",
INIT_24 => X"FFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFFFFFFFFFFFFF552A974",
INIT_25 => X"0010000000000000000000000000000000000000000000000007FFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0804154BAF7FFFFFFFF",
INIT_2B => X"FFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA",
INIT_2C => X"00007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000AAA2FFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804000100000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A",
INIT_31 => X"04174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAF7FFFFFFFFFF",
INIT_32 => X"FFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E974AA08",
INIT_33 => X"AAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA2FFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"5886C0201A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"0005EE040057700F40D08078500000D9218020407F0000BB8018A2FC380BEAC2",
INIT_05 => X"F0F817FFFE400800020224000405F7FFE0124002FFE1E0C517FF09111212F300",
INIT_06 => X"400000409120338860900482404FFFFC000000001FFC0832050E00047F97870B",
INIT_07 => X"00246801C41C3E81E872C8FFE900FC31348EFDF03BE15E22DA07FF92C2041020",
INIT_08 => X"6220280D2B025988311AB14155421006891A1089F6E200000022C140068EB902",
INIT_09 => X"0002021FFEFBC80000000077FF184B03010004002FE1F2900201000000FFDFFF",
INIT_0A => X"0006FFEA002020626995FBE077430001E7320006F87D7FA84024B0225A890FFF",
INIT_0B => X"241C482B20400CC52492710CC80060020A81BFE41FF0C2060481200180000000",
INIT_0C => X"040430404304043040430404304021820218210018C24110A860006C620C0312",
INIT_0D => X"001002001804800000952800001FFBF040C088669070510C90C1430404304043",
INIT_0E => X"1FFEAFFF805025E00853B92588000400020001000020A8018008002000014030",
INIT_0F => X"148484054395E27E428002A4200397E07E422002A420100382FCC30832A16382",
INIT_10 => X"788417000397E07E428002A4200395E27E422002A420110A51C01C0590401486",
INIT_11 => X"1A2490040590C08120558C1759BE1C05A0400383808800DA1929F728641100C0",
INIT_12 => X"00136006000215EA0A4833A32C8832050028603050014031B3950000C90A51C0",
INIT_13 => X"658280009A2030108B14AC05C00112405222088B8332C140004D101800CE7200",
INIT_14 => X"B6808060201281004228996085F10020180C030880D11019CE4000026C00C006",
INIT_15 => X"49DC7143F01C04240030720641E0A028996483A17204680410A04104A2659196",
INIT_16 => X"1000080080000000000002001201F7FFC0011C2F81A48080CA32800A0108152A",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"0000000000000000000040100401004010040100401004010040100401004010",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080002010FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA08",
INIT_33 => X"F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"0000745C200801000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"0001E6000053300F00D0007810042140C00000407F0000BB800000DC3801EA00",
INIT_05 => X"F0F8033FFE000000000000000001F17FE01240009BE1E00003BF00000000F300",
INIT_06 => X"000000009120110020100002404FFFFC000000001FFC0000010E00007F878701",
INIT_07 => X"00102050840950002802C87FC800FCAA035400001B918600C207FF8000000000",
INIT_08 => X"6234AD280B02500063AC2840001610020408178B600C24000136496087300042",
INIT_09 => X"00000007FEFBC00000000077FF000B00000000002FE0000000000000000FDFFF",
INIT_0A => X"0006FFE80000015406A800003388000025000002387D7F804024B0224A8107FF",
INIT_0B => X"20502000200000400490510CC00040020201BF441FF0C0000000000180000000",
INIT_0C => X"040030400304003040030400304001820018210018C0411020600048620C0300",
INIT_0D => X"800B00000000000000000000001FFBE0008080641060400C00C0030400304003",
INIT_0E => X"1FFEADFF80002080000000208800000000000000000020018000000000000004",
INIT_0F => X"009181008024A00043601100210024A00043C0110020901382CCCB28B0806202",
INIT_10 => X"040A03080024A00043601100210024A00043C01100209240C840C201D0210840",
INIT_11 => X"A604E0080820009908008341B000A8212070082002890010068320860C920180",
INIT_12 => X"00800082041205EC00044C1ACB66C37542082030281E0580001012811A40C840",
INIT_13 => X"27A004300004103160DB3005E000618040C022000593D002180002090166B406",
INIT_14 => X"FF20406040084210C062000C2A2DDD00180C04504086002CD680C0100010480B",
INIT_15 => X"04295C98F80400008040CC0582169022000C2876C404780028500160880012BB",
INIT_16 => X"0000000000000000000000000001F7FFC001B823018F00880008805241060208",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9EF9EFB263CC3090CABAEBAFF96857757B73E6089966B9EF9D5A220CC8000000",
INIT_1B => X"0F0783C1E0F0783C1EFBEFBEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF",
INIT_1C => X"0000783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2010000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020100000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA00",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00004000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"4909E6093253306F82D0007C80000000080E01007F8020BBC00040DC3801EA00",
INIT_05 => X"F0F8033FFF0240012C1400080291F17FF01241009BE1E00203BF80800000F392",
INIT_06 => X"0DC00CC0992033A062116E82404FFFFC0E0801101FFC0000010E08A07FC78701",
INIT_07 => X"00000000000000002802C87FC800F8000000000019810600C207FFF3C410D841",
INIT_08 => X"E8002000080281000008A0000014100200081000000000080480AE0000002000",
INIT_09 => X"80040007FEFBE031018C31F7FFBAEBC0020008086FE0000100280800000FDFFF",
INIT_0A => X"0006FFF800C04000000000003300800005000032387D7FE94FBEF2B2CB8DA7FF",
INIT_0B => X"20100000200000400490D10EC00040220201BF441FF0C0600000000180000000",
INIT_0C => X"04003040030400304003040030400182001821001DCCC31222730A49620C0300",
INIT_0D => X"000000000000000000012800001FFBE0008080641062400C00C0030400304003",
INIT_0E => X"1FFEADFF805025C0304001E58906088304418222C108A009A090400000000000",
INIT_0F => X"00100100000480000200100000000480000200100000100380F0C30830A06302",
INIT_10 => X"0008000000048000020010000000048000020010000000004040000010000000",
INIT_11 => X"0004000000000008080000011000000020000000020000000001200000100000",
INIT_12 => X"000000800002018C010000020800000800122000000004004000008000004040",
INIT_13 => X"2080000000040000001020020000000000800200001040000000020000021000",
INIT_14 => X"1000008001000000800200000021000020100000000200004200000000100000",
INIT_15 => X"0008400000000605000000000200000200000020400000000000002008000002",
INIT_16 => X"226410410346010000000400A011F7FFE0031823010400800000800001840000",
INIT_17 => X"2088220882208822088220882208822088220882208822088220882208822288",
INIT_18 => X"0882208822088220882208822088220882208822088220882208822088220882",
INIT_19 => X"17FFFFFFFFFFFFFFFFE088220882208822088220882208822088220882208822",
INIT_1A => X"0492410A048029890AD34D35FDD144A50CB5462D14997BE09E760AED04040000",
INIT_1B => X"6231188C46231188C49249249249249249249249241041041041041041049241",
INIT_1C => X"000B158AC562B158AC562B158AC562B158AC562B158AC562B158AC562B1588C4",
INIT_1D => X"0000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"94A7B2B1450000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"6FEBEF5FEC737AFBC6F85FDEB220109E1FEFFFE3FBA7FDFB9BD301DC3FF5F0D2",
INIT_05 => X"F0FFEB3EFFF7FDED3FBFF6A84383F177F5FB7FF59BE1FF980BBBB7FE6D21F3DB",
INIT_06 => X"FBE564C71268F3BBF5FBFC2A427FFF7C3E3A74667FDDB7FB870FF30FFDEF87F5",
INIT_07 => X"3BC18306396FBEC14489737FDC00B13BB79DFDB83BF4112AF205FFBDD3AFB93A",
INIT_08 => X"21E4391909B381B0B1F8E041051831FA3068D77E000030021324620C0B9C2060",
INIT_09 => X"D13D980FBEFBEBF30B8D79FF7F451F33CFD60FE8FFFDF54003B1D4223B4FFDFF",
INIT_0A => X"B5AFF7CFACFAFE776F39FF7077E29D83CFAB300B017F5FFE6FBEF73BEFB967FB",
INIT_0B => X"737AF3FD62601EDC25B3533DCEB07F262213FFC67FF1C7FBFB5EC9478D5DA3A3",
INIT_0C => X"5E3035E3035E3035E3035E3035E981AF181AE315BDDCC3B336F7C548667D47B7",
INIT_0D => X"100C0E60FB9FC3A80EF69A004DFFFF7FF5F9A06E19F4DA0E80E903DE3035E303",
INIT_0E => X"7FFFF9FF8FAFAA3ADEBFB9726BAF5FD7AFEBD7F7EFFD7ACDB7F947F0EA035CF6",
INIT_0F => X"0080A40403E8BD8002000FC02003E8BD8002000FC02010979AFFE36C36B86702",
INIT_10 => X"EE00034003E8BD8002000FC02003E8BD8002000FC020037B0040A00010003E02",
INIT_11 => X"C00400003D80008160400FD81341C00020003B80008C00801EF0285380100000",
INIT_12 => X"81038406809677FA080468C46A81080581002000780C8001C8100201037B0040",
INIT_13 => X"90D162001C803411FC0024080001F80040026C0807C868B1000E401A01F11909",
INIT_14 => X"10503A00003E020042AC080CEB01228A80000F600080123E232130407080D00F",
INIT_15 => X"7520750001064180807868000110C02C080CFA0042400000F8800105B02013F8",
INIT_16 => X"FF7EFEEFF3EEC3FF7FBFFBCB7FFFFEFFE00BFF7FEBF420800EC0CBEE61F81008",
INIT_17 => X"F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F7FD",
INIT_18 => X"5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7",
INIT_19 => X"37FFFFFFFFFFFFFFFFF5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F",
INIT_1A => X"A61861BAF15EAA6AFC38E38EA3AD8ADE7A48F0B366429F434AA9FC376DAE4432",
INIT_1B => X"130984C26130984C261861861861861861861861861861861861861861869A69",
INIT_1C => X"0000984C26130984C26130984C26130984C26130984C26130984C26130984C26",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"1085B0B041000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"6FAB975B6470BAF386C87A9CB00000001FEF9F23E3A7BDE79B5101D23FB5C0C2",
INIT_05 => X"C8FFCB38FF35B44C25ADE72041A3F147F5FB7F759B91FB880BA3B6FE2921CBDB",
INIT_06 => X"B98420C71408D113956AFD0842FFFC7C3032646EFF1DB7FA868FE30EF1CE47E5",
INIT_07 => X"0041830600640C415004637FC4003021259CFDB01BF80028E001FF8251AB9D1A",
INIT_08 => X"200822020842203000082050000110023068D030000028200000008400000051",
INIT_09 => X"90A4880E3DF7E2FB0B8E717C7F411F3BC6D60B60FFDDE440018AC4AA3B0FD1FF",
INIT_0A => X"042787C5AC5ADC424B39FB6073D00D8048A31008017C1F826FFEF41FEEB027E3",
INIT_0B => X"7BEAF1C152201A4C05B7531D56B05B06A213FF863FF5D5F9FB5E8847A0702606",
INIT_0C => X"0D1030D1030D1030D1030D1030F0818688186B51BFDCC39732F3554866AD57C3",
INIT_0D => X"10080A20ED1D41880CC61A0044DFFC6EB5BCA06F18FC5A0E00F0038D1030D103",
INIT_0E => X"3FFE91FF98AEAA1AC6AC9A3A4AAD5B56ADAB56D5AFD572C597B147506203E8FC",
INIT_0F => X"0000260403C8948002000EC0000BC8948002000EC00010878AC3CB8AB8857202",
INIT_10 => X"EE0000400BC8948002000EC0000BC8948002000EC000097B0040200010003E02",
INIT_11 => X"400400003D80000070400DD81041400020003B80000410801AF0204180100000",
INIT_12 => X"010384008086378A080428C46A80080081002000780C800188000301017B0040",
INIT_13 => X"909042001C800409FC0020080001F80000007C0807484821000E400205D11101",
INIT_14 => X"10100A00003E020000BC0808EB01020280000F60000002BA222020407080102E",
INIT_15 => X"7520750000024080807868000100403C0808FA0040400000F8800001F02003F8",
INIT_16 => X"EF3AF6AF6389C2FE128971AB2DDDF8FFE0031B776BF4208006C0C92621F81000",
INIT_17 => X"D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B5",
INIT_18 => X"5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56",
INIT_19 => X"3FFFFFFFFFFFFFFFFFD5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D",
INIT_1A => X"0000001E0080397908000000A48710B4080240E543021B438A010825238B443A",
INIT_1B => X"4020100804020100800000000000000000000000000000000000000008200000",
INIT_1C => X"000A05028140A05028140A05028140A05028140A05028140A05028140A050080",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"8C2100804900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"02000100440408002408008002221000204116A280000F000001400000100010",
INIT_05 => X"00000000001265050080C000190002000000005C0000000A0000002C20600000",
INIT_06 => X"14016012000C405280200008001000011110012220009A88800009A880000000",
INIT_07 => X"0048912242288100800102000400010208000000040000082000002400814008",
INIT_08 => X"0A010040401080308400821155540001122448142491008A0049120408402210",
INIT_09 => X"04080A000000124058200408000880004440004080160C4100A8580099400000",
INIT_0A => X"4A50000080080E041000000008000C81000110010500002000000180001C8000",
INIT_0B => X"110091500020B408810000100200020408B0000020000081B2C208420ADA5353",
INIT_0C => X"5814058140581405814058140580A02C0A02C004800210C19808400500010009",
INIT_0D => X"10040860B188C0A80653020005A004039010280000800B00100040D814058140",
INIT_0E => X"600010000280000802050010660001000080004004900204020105302A000C42",
INIT_0F => X"0000A00000081480000001400000081480000001400000800C01082082210500",
INIT_10 => X"0000024000081480000001400000081480000001400000010000200000000000",
INIT_11 => X"4000000000000001400000080041400000000000000C00000010004180000000",
INIT_12 => X"0100000480802A40000000400000080081000000000000004800000000010000",
INIT_13 => X"1010420000002400040000080000000000024400000808210000001200010101",
INIT_14 => X"00100A0000000000028400004000020280000000000012002020204000009000",
INIT_15 => X"1000000000024080000000000010400400004000004000000000000510000040",
INIT_16 => X"8408420430E699AA42A1508104EA08000000810020000000044001AC20500000",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_19 => X"8000000000000000000010040100401004010040100401004010040100401004",
INIT_1A => X"20820800D41A8283AC618618EF1088160885001234B96061CCDEC4D205061170",
INIT_1B => X"6030180C06030180C08208208208208208208208208208208208208208208208",
INIT_1C => X"000B0582C160B0582C160B0582C160B0582C160B0582C160B0582C160B0580C0",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0803B2814D0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"26E1E905CC574828C4F85FC600000016004F77E2F887CDB80BC340DC07D1F000",
INIT_05 => X"F007E33E01D26CE43A92F2880B01F37011E93ED49BE01F1A03B8972E6D20F049",
INIT_06 => X"5AA06002026872BAE0B1282A005FFF001E1870223FC3BFC98101F109FC6780F1",
INIT_07 => X"3BC081023B233E804488527FDC008019968D74982C94110AF204001BC285A828",
INIT_08 => X"01E4191901A101B031F84000000831FA1028575A000110800124600C039C0020",
INIT_09 => X"C1111A0782082B50080508FF00048B124D4005C8AFF4154102914800110FFC00",
INIT_0A => X"B5AAF00A80A82C332D18ED301D229C82C7A93002017F405C409A42A9A51547F8",
INIT_0B => X"1158936D20601A98A10200308A002E240010BFC0600002AFFBE249420555A2A2",
INIT_0C => X"1A3401A3401A3401A3401A3401A9A00D1A00C000850400A11414C005005000B5",
INIT_0D => X"10080C60AB0F42A8046282000DBFFF13D059280201948B029029409A3401A340",
INIT_0E => X"6FFFF8000F8F80281A16A1504302058102C0816244B82A0CA25907D0AA015874",
INIT_0F => X"0080A40000283D80000001402000283D80000001402010901A7D694494192200",
INIT_10 => X"0000034000283D80000001402000283D80000001402002010000A00000000000",
INIT_11 => X"C000000000000081600002080341C00000000000008C00000410085380000000",
INIT_12 => X"81000006809076B2000040400001080581000000000000004810020002010000",
INIT_13 => X"1051620000003410040004080000000040026C00008828B10000001A00210909",
INIT_14 => X"00503A000000000042AC00044000228A8000000000801204212130400000D001",
INIT_15 => X"1000000001064180000000000010C02C000440000240000000000105B0001040",
INIT_16 => X"964C4A44A0C689FF3F9FFEC5D6DBFE0020096528A0B000000CC043EC60780008",
INIT_17 => X"6058160581605816058160581605816058160581605816058160581605816258",
INIT_18 => X"0581605816058160581605816058160581605816058160581605816058160581",
INIT_19 => X"17FFFFFFFFFFFFFFFFE058160581605816058160581605816058160581605816",
INIT_1A => X"AEBAEBFFF7FEFCFDF7FFFFFF5DE7CFCB773FFEFBFF3C7E1E779FFEFFF5060030",
INIT_1B => X"F7FBFDFEFF7FBFDFEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEB",
INIT_1C => X"000FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEF",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9E79E7BAF7DEBAFAFEFBEFBFFBFFDFFF7FCFF0FBFFDFF7EFDDFFFEFFE8000000",
INIT_1B => X"7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"0003F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"1084B030000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"6DA986092050306382C05A1C900000001FAE89016387B2A38B5000D03FA1C0C2",
INIT_05 => X"C0FFC338FF008048240426200081F147F1FB7F289B81FB8003A396D20940C3DB",
INIT_06 => X"098000C51000910100006C00426FFC7C202060445F1F2572060FE82671C607E1",
INIT_07 => X"0001020400440C41C000617FC0003021259CFDB01BF00020C001FF8040009800",
INIT_08 => X"2000200008020000000820440000100220489020000020000000000000000044",
INIT_09 => X"8004800E3CF3E0B1118C31747F000B33820209206FC9E80000000000220FD1FF",
INIT_0A => X"000687C0044040424B39FB6073C0010048A20000047C1F804FBEF01BEE8027E3",
INIT_0B => X"204A608142002A440492530C401049020221BF861FF0C06C493C800580000000",
INIT_0C => X"04003040030400304003040030600182001821011DCCC31222730048620C4382",
INIT_0D => X"000802004815010008840800405FF864008880661874500E00E0030400304003",
INIT_0E => X"1FFE81FF880EA000400098200C04080204010200810020C180904240400340B4",
INIT_0F => X"0000040403C0800002000E800003C0800002000E8000100780C2C30830806202",
INIT_10 => X"EE00000003C0800002000E800003C0800002000E8000017A0040000010003E02",
INIT_11 => X"000400003D80000020400DD01000000020003B80000000801AE0200000100000",
INIT_12 => X"000384000006118A080428846A80000000002000780C800180000201017A0040",
INIT_13 => X"808000001C800001F80020000001F8000000280807404000000E400001D01000",
INIT_14 => X"10000000003E020000280808AB01000000000F600000003A020000007080000E",
INIT_15 => X"652075000000000080786800010000280808BA0040000000F8800000A02003B8",
INIT_16 => X"223010010308025410082404A015F0FFE003182701B420800280C80201A81000",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_19 => X"17FFFFFFFFFFFFFFFFC080200802008020080200802008020080200802008020",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000080040",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"88280C4C7B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"00160090920C04800904848262220277E05152B280780D407428E723C01E1400",
INIT_05 => X"0F001CC000890026105810941C5C06800E008057641E00473C40680D32330C00",
INIT_06 => X"82541A028D584E40CB0583CCA0100000161F84322000DA8C40F003C80030780E",
INIT_07 => X"BF70E1C3BBBB1138AF7F888025340C0888430047040FEE182CA00044BC5827C5",
INIT_08 => X"CAFC1F1F07F0FE1C94F65B11555EAFFC1C306758B24197ABCDA467F2C9CF9B32",
INIT_09 => X"4FFB4730000011420A61080800B6E0C464258094101606D5A47A2A2098B02000",
INIT_0A => X"446000304A0488111084048E082D0ED020119D35F900002FB00105C01036D800",
INIT_0B => X"1FA599581D3A9583C105A892112C04C0A898403120071501A6C32222068A3050",
INIT_0C => X"789E07A9E0789E07A9E0789E070CF0184F038850A21008E514845AB510D0106D",
INIT_0D => X"9A95E954868AD0E52273F4AC2180000808061C01C48B0F81380CE0F89E07A9E0",
INIT_0E => X"4001120055704FC4A1624487E2489024481224091282C4300942A19439481842",
INIT_0F => X"5D65C3E3F01F52FFC1E0013C1F801F52FFC1E0013C1F8090423D38A18E3B15C9",
INIT_10 => X"118796BE001F567FC1E0013C1F801F567FC1E0013C1F9085DFBF7E15C06101C5",
INIT_11 => X"7E30F00C0270F3751F1FD00FECBF7E25C0700463E17B2C7F811FD7ADECC381C0",
INIT_12 => X"4190626D6491063597F9177B956EF378D33E4030061341F077C571F8F885DFBF",
INIT_13 => X"7F328E3082636B2807FFD80FE00007E03F7207D3E03F9167184131B5C40FE647",
INIT_14 => X"EFA0CAE06101C53E3647D3F144FCDD22B81C0098E57D9081FCE8C8520C4DAE20",
INIT_15 => X"1ADF08DBF81846A540049707E0FE3307D3F141FFB45478040570EED41F4FE047",
INIT_16 => X"C189601208A1502B4AA5584B4068000019A80098120BCA4C617635C938574FF3",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"A800000000000000000902409024090240902409024090240902409024090240",
INIT_1A => X"08208208831042720EE38E38AAF9C4C704DAB63A6D58B3C10BAE8E789AA09424",
INIT_1B => X"7C3E1F0F87C3E1F0F82082082082082082082082082082082082082082082082",
INIT_1C => X"0003E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F8",
INIT_1D => X"0000000000000000000000000000000030F007FFFFFFFFFFFFFFFFFFFFFFF900",
INIT_1E => X"155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AEBDEBA0000000000000",
INIT_1F => X"7FD5545FF8000155087FC0155F7D168B55007BFDF45085168ABA002E82145085",
INIT_20 => X"55568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D7FFFE1000554214555",
INIT_21 => X"FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF7FFC00100800175555",
INIT_22 => X"0002E974BA5D5168A00A2D142155005142010FFAE820AAFF842AABAA2AE95545",
INIT_23 => X"AAFF803FFFF5D2A821550000000BA007FD55FF5D7FC0145007FD740055041541",
INIT_24 => X"FFF082EBDF455D5142000082E82145FFD17DFEFFFD168BFFF780000BA007FE8A",
INIT_25 => X"FE3F000000000000000000000000000000000000000000000AAFBEAA00007BFD",
INIT_26 => X"6F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEBDFD75D2AA8A80EA8E2",
INIT_27 => X"1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B68B551475FAF6D1C55",
INIT_28 => X"7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA0000542A0070071C50BAFEF",
INIT_29 => X"B8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A8010E004924874825D",
INIT_2A => X"EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0120155EA568E870BAE",
INIT_2B => X"7ABA497A82FFAFD2A82485FD2415A105C21451ED42A002545E055FFBE81D0BE8",
INIT_2C => X"00B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6A5C7E3DFFFE90B45B4",
INIT_2D => X"F45592E88A0AFE80A8B0A0000000000000000000000000000000000000000000",
INIT_2E => X"A1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE975EFAAAAB5E1AF3AABF",
INIT_2F => X"1CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB65F520EBE9EF67D7BE",
INIT_30 => X"034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EBC11472800752117082",
INIT_31 => X"968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F3142341D5DEEBEF55080",
INIT_32 => X"7D58AC448B69C30E02116220415A9540AA854140A0A2047F353AAF6C77F7F20D",
INIT_33 => X"56EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7C91565455C141E4188",
INIT_34 => X"F0000001FF0000001FF01EABC4B8014174FF7DA80F52FEDE6BE93172D7D625B5",
INIT_35 => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F",
INIT_36 => X"0000000000000000000000000000000000001FF0000001FF0000001FF0000001",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000100000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"CA1800080848B0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000010822C00803804000001999EF9C00040B0002000001000640200001018",
INIT_05 => X"08000000000100030008010468220A0004000000001000032000200002100800",
INIT_06 => X"8201961000060444010081002080000080820100000008004880000000284000",
INIT_07 => X"210C18306788C0089409800001140082000100010405000410A0000010082500",
INIT_08 => X"0A48903121780004C6000311555521F183060AC564BF818B5EDFDE0044600301",
INIT_09 => X"45B103200000140802234800000584000004808400020011A4581A2200002000",
INIT_0A => X"021000000800810400000402083000510000050020820036200005C00026C000",
INIT_0B => X"40000002000A008182200000002404400000000000010500008020A022220040",
INIT_0C => X"68064680646A0646A06468064690321503234204020018200404010784700404",
INIT_0D => X"C417C16004C0B838221090240180000801000C8800000190191064620646A064",
INIT_0E => X"6000000010200200802100022008100408020401020040100142200E0E08A20B",
INIT_0F => X"0021E300B000000781E00140018000000781E00140018000002430E30E0615C9",
INIT_10 => X"0000024E0000000781E00140018000000781E0014001908400005E11C0610000",
INIT_11 => X"3C30F00C000000155800D00000003E21C0700000000F00118000000468C381C0",
INIT_12 => X"40900004A400081401A0000004041218503E4030060000004804318008840000",
INIT_13 => X"01208C30800025200003D807E000000000725201600090461840001340002606",
INIT_14 => X"0F00C0E06100000012D2005100409520381C00000005920004C0C81200009A00",
INIT_15 => X"00120850B8180625400400000010711200510004B41478040000005548016000",
INIT_16 => X"40002002080000000804000A0000000011A000100208C008611430A000040250",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"0800000000000000000100401004010040100401004010040100401004010040",
INIT_1A => X"8A28A2AC8090C69606492492C09945235D5F7E2A5040B80E1C863A2958000500",
INIT_1B => X"DD6EB75BADD6EB75BAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A2",
INIT_1C => X"0002E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BA",
INIT_1D => X"00000000000000000000000000000000C0FFFFFFFFFFFFFFFFFFFFFFFFFFFC00",
INIT_1E => X"FE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5555550000000000000",
INIT_1F => X"D1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7AEBDF455D2EAABEFF7F",
INIT_20 => X"5000015500557DF45AAD1400BAA2AE801550051555EFF7AA95400552AAAABAFF",
INIT_21 => X"F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB5500517DF555D2EAAA105",
INIT_22 => X"5552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBAFFD540155557FD5400",
INIT_23 => X"10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAABAFF842ABEF5D517DF5",
INIT_24 => X"E105D2E954BAF7AE80010082A97410557FEABFFAAFBE8BEFAAD1575EF557FFFE",
INIT_25 => X"056A0000000000000000000000000000000000000000000005D7FFDF4500043F",
INIT_26 => X"BDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC51C7A2FBD5490BFD1C",
INIT_27 => X"4924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA974BAF7FFEFB45FFAA",
INIT_28 => X"DB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2080BEF495FC71D5412",
INIT_29 => X"FD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4002D082082AB8B6DBE",
INIT_2A => X"487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF78E021FF1471FDEAAF",
INIT_2B => X"FF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545A2DA3FB7DAAD4AAAAF",
INIT_2C => X"00547AB8F550A8010E00492487482FFFE82A85EBAE2FFC55554ADBD7A2FFC7BE",
INIT_2D => X"545AAFBF7400FBF9424F70000000000000000000000000000000000000000000",
INIT_2E => X"74AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E5400021EF005162BEF047FD5",
INIT_2F => X"225FF5843404547184164AA5D2EBEEB0A2D555410D3555714F8338AAAA1D0AE9",
INIT_30 => X"409000512AEABFFDF79DCBF755962010BDCBBC21455D7FEABEF75550ACBB7582",
INIT_31 => X"0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3FFEAAEB083BC1000FF8",
INIT_32 => X"BD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF801F8BA0C57740BDAA",
INIT_33 => X"DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF5D16BABAA3EBC3157A",
INIT_34 => X"0000000000000000000596EBEF55080034E0A592A4AD00FB863550229BCABEB7",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000100000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0812",
INIT_01 => X"A145A00810790848048044A54E404340404000720885800802000906E4910200",
INIT_02 => X"5C010802020408040C455850AA055254090541A111200A104A0000000908B510",
INIT_03 => X"182002200C00004485264A001214912803150020218808002440854288890550",
INIT_04 => X"210302048014100160806B08702010102722C9E0412200651102418214049492",
INIT_05 => X"88510910540008812C06010018204342A58A08011290A1120A81230240018DCA",
INIT_06 => X"47450000022480090000210002A54C282122040CC9082D530085224410AA4204",
INIT_07 => X"2101020423408900940C402A900011012D41D518044C10025000AA8A50043D00",
INIT_08 => X"214912534123010085008010141521F020409260000100A00004428808102010",
INIT_09 => X"519D12041551589141A539C42A4C9608080004801700D10100311820A848E0AA",
INIT_0A => X"0244C28C000002025A81AE3048321002A700200900160AE42CAA839AA90442C1",
INIT_0B => X"42300225604004D080251121D0000400880178044355940A498C400004A00545",
INIT_0C => X"4F240472404F240472404D240441200692022B41365E53340EC6940564D012D6",
INIT_0D => X"00000620500403080A919000038AD03001C5080D1108C1009001404524045240",
INIT_0E => X"02AA40AA902408000010002220040C000201030201200C818098402082020438",
INIT_0F => X"0080A0000140000002000140200A8000000200014020100280E469C698353000",
INIT_10 => X"000003400A800000020001402009400000020001402008700000000010000000",
INIT_11 => X"0004000000000081400004C00000000020000000008C000010A0000000100000",
INIT_12 => X"0000000680004188000400840080000000002000000000004810000001420000",
INIT_13 => X"0000000000003409280000000000000040025000030000000000001A05100000",
INIT_14 => X"000000000000000042900000A100000000000000008012A2000000000000D026",
INIT_15 => X"4420300000000000000000000010C010000098000000000000000105400002A0",
INIT_16 => X"126000808200505448342228120090554000E00000000000088000A000000000",
INIT_17 => X"004010040300C0300C0300C0100401004010040300C0300C0300C01004010240",
INIT_18 => X"0400004000040000C0200C0200C0200400004000040300C0300C0300C0100401",
INIT_19 => X"9FC0FC0FC1F81F81F800C0200C0200C0200400004000040000C0200C0200C020",
INIT_1A => X"0410411823A4301040B2CB2CBACB002009C6B860185AA1491B0E2863E8001100",
INIT_1B => X"4A25128944A25128941041041041041041041041041041041041041041041041",
INIT_1C => X"03F25128944A25128944A25128944A25128944A25128944A25128944A2512894",
INIT_1D => X"00000000000000000000000000000000F0F007FFFFFFFFFFFFFFFFFFFFFFFC07",
INIT_1E => X"415410AA8415555087BFFF55A2AA800BAFFAE9540008002AA000000000000000",
INIT_1F => X"FBEAABA5D7FE8B555551421455D0002145552EBFEBA007FC21EFA2FFD75EFAA8",
INIT_20 => X"2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F784155EFA2AEBDEAAA2",
INIT_21 => X"5D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BAA",
INIT_22 => X"55D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AAAAAAAAAAAFFD157410",
INIT_23 => X"FFA2D17DFEFF7800215500557DF55AA80001FFAA80001550055575EFFF840215",
INIT_24 => X"0AA082EAAB5500517DF555D042AA10A284154005D0015410085568A00FF80175",
INIT_25 => X"8A2A0000000000000000000000000000000000000000000005D00020AAAA8002",
INIT_26 => X"C51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA800AAFFAA9543A08003",
INIT_27 => X"0105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF49040017D5D20B8EAA007F",
INIT_28 => X"A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492AA8BC7EBDFEAFEFFD0",
INIT_29 => X"6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6FFEFB6D555578F7DB6",
INIT_2A => X"0155C51D0092A071555D5E3AE821D00001FF0871C016DBED1FDE90E3A497492B",
INIT_2B => X"8007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6DBE8F401D7B6A000147",
INIT_2C => X"00410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C5BE8555400550A3842",
INIT_2D => X"0AAF7AA954AA00042AAA20000000000000000000000000000000000000000000",
INIT_2E => X"21EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE975EF005560B55F7AA80",
INIT_2F => X"A8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BEABEF057D68F5F5A000",
INIT_30 => X"BFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D57DF55D7AABFF5428AC",
INIT_31 => X"D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002CA8AA80800020AAF7F",
INIT_32 => X"680800FFF7AAA155F595542455512A975455D3AA8A005500151FF0C57401E5F3",
INIT_33 => X"7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A2AA801455D7FE8BFFF",
INIT_34 => X"00000000000000000000C3BC1000FF8409000512AEABFF5D79FCAF774AE005BE",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000200000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380206",
INIT_01 => X"014C9A40408001683C0462C99E004B61404040028804A0080A000D16A0990A0C",
INIT_02 => X"4809A902031800444460589C66E331352180D468B8240E600C0081110B80ACD0",
INIT_03 => X"DA14C2210C0001D235834A0648D60528330006810A80881068A80C029CC56330",
INIT_04 => X"20886819A02740ECD2107364B37569100A04C1E01CA52010990240420E205A08",
INIT_05 => X"5831803532410000260E272058232259954369000A506912018CA582480038D1",
INIT_06 => X"8381A014000200AC2190ED0002ACD99881822144C5A409430682800046294140",
INIT_07 => X"218408142740E2C0948C3066500071913209CC8004640102D003999552083D20",
INIT_08 => X"00409231296AA180C2000110001521F0810A92E7402F00AB0016CA080C600111",
INIT_09 => X"41B112014D30E43802A76DD09905882B010605A01A4941010211088A2A43A399",
INIT_0A => X"4A12D9820880832264119D004860900104002008000F399606BC07998BA546AC",
INIT_0B => X"42522013604080D084A01001C8302D00008153000731C3000988C0040A224110",
INIT_0C => X"602406824068240602406224068920151203030032545B7404D7804566594796",
INIT_0D => X"080600E04C442068088590000999C8E84041086C001091009001406824060240",
INIT_0E => X"E6660599902600209021204A010E1C850C428521C208480021D842081A03E231",
INIT_0F => X"0090000003200000000010002008A00000000010002008038666928B28A65300",
INIT_10 => X"000801000A200000000010002009E0000000001000200A380000000000000000",
INIT_11 => X"0000000000000088000002D00000000000000000028010001620000000000000",
INIT_12 => X"0000008201021C88000048800280000000000000000004000010000003600000",
INIT_13 => X"8000000000041019980000000000000040802000068000000000020805B00000",
INIT_14 => X"0000000000000000C020000C8300000000000000008200AE000000000010402B",
INIT_15 => X"41003100000000000000000002008020000C3800000000000000012080001298",
INIT_16 => X"737420C20A01405468360022201185CCE0128410820000008088021C40A00008",
INIT_17 => X"2108721085218852188521885218852188521887210872108721087210872308",
INIT_18 => X"1086214872108621C852188421C852188421C852188721087210872108721087",
INIT_19 => X"26AA555AAB554AAB5561C852188421C852188421C85218842148721086214872",
INIT_1A => X"0410412881D0B0000092492480A981E063C638321450A08899A62C314A810508",
INIT_1B => X"EA753A9D4EA753A9D49249249249249249249249249249249249249241041041",
INIT_1C => X"BC4351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A9D4",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF82A",
INIT_1E => X"02AA00AA843DF55FFAA955EFA2D168B55557BEAA000055420000000000000000",
INIT_1F => X"5568A00087BE8BFFA2D155410AA8415555087BFFF55A2AA800BAFFAE95545080",
INIT_20 => X"D0002145552ABFEBA007FC21EF007FD75FFAA841541008002AB55AAAA955EF00",
INIT_21 => X"5D7FC0155005168B455D042AB45F7FFD741000042AA10AAAABFF5508003FF555",
INIT_22 => X"A5D7FC2010A2D1575FFF7AA975555D2E80145F78415545082EBDEAAA2FBEAABA",
INIT_23 => X"FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABFFF7FBEAB55F7AABDEB",
INIT_24 => X"B5555557DF55A2AEBDF555D2E954BA002EAAABA002A821EF5555554AA087BC01",
INIT_25 => X"203A000000000000000000000000000000000000000000000082E820BAA2FBEA",
INIT_26 => X"800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6FB7D5D7FEAA3808554",
INIT_27 => X"E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E1557D1475FAF45BEAA",
INIT_28 => X"AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2FBD55D7BE80004AA1E8",
INIT_29 => X"C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FFF5D0438140E2FA38B6",
INIT_2A => X"EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75D0A901FFFF801557D1",
INIT_2B => X"74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB455D20BDE00EBAAA8BC7",
INIT_2C => X"001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125FF002EADA921420871D",
INIT_2D => X"FFF5D7FEAABA0051400A20000000000000000000000000000000000000000000",
INIT_2E => X"75EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAAB55A28408145AAFFFF",
INIT_2F => X"D7145FBB8020A35D2ABEF55F7800015F087FEAA00007FEAB55FAD568AA2AFAE9",
INIT_30 => X"5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF55042AAAA007FD55558A7B",
INIT_31 => X"040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057968F575D003FF55F7D",
INIT_32 => X"52A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AAFFD5145FBAC9755F05",
INIT_33 => X"052ABFE10550415557085540000005156155FE90A8F5C082E974AAF7D57DF455",
INIT_34 => X"00000000000000000005500020AAF7FBFFFEF04552ABFFFF843FFE77C80825BC",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000100000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804002061080A284201081034809800A00230340007833522C82D04A16002",
INIT_01 => X"80439982183828490400050E12000340403008418984014902030106A0D10204",
INIT_02 => X"480108A000000000446418E01E80F00A41043118680402000800000009882390",
INIT_03 => X"0CA080210C0000408006480002001120260012603000000030808900888100F0",
INIT_04 => X"4403A609A055306B82C0705800CEE510082AC0A16B0350E3808041D03865D002",
INIT_05 => X"C0F20B36F0000901240626200820E26780E244A19A41E4020BAB06404001D312",
INIT_06 => X"434420151220118900806922406C3C7800201448DD9D2870020F228075A60715",
INIT_07 => X"2181000023480040840C001E180030032009700024641002C00187A440047C00",
INIT_08 => X"084830110160208004000001101121F220000260000100AA0004408000000001",
INIT_09 => X"519102063DF3E02B100B097407448F200A0209A041CA290102130C8800466478",
INIT_0A => X"8543D048006040064010E4007F62110105002002044007846124E0A00E0DC1EB",
INIT_0B => X"60020291404024808030512C40106D022203B1445810856A019400058F8404B5",
INIT_0C => X"052430D24305243052430D24304121A6921863013FD8807626EE000D64540284",
INIT_0D => X"28081080508104400A00800009B878680000880C1160410C90C143152430D243",
INIT_0E => X"81E0E18790012A00080102280800000202010102810020018098404110020004",
INIT_0F => X"0090000005E0200000001000200C6020000000100020000390E6C30830806204",
INIT_10 => X"000801000D20200000001000200EE0200000001000200A6A2000800000000000",
INIT_11 => X"8000000000000088000003B00100000000000000028000002EA0001000000000",
INIT_12 => X"80000082000251D80000C0044280000100000000000004000010000003282000",
INIT_13 => X"00002000000410121800040000000000408030000B8000100000020806F00000",
INIT_14 => X"0000100000000000C030000C9000008000000000008200FC000010000010403B",
INIT_15 => X"A500100000000100000000000200803000042E000200000000000120C0001590",
INIT_16 => X"30000800002400044934040AA231B63C20530801000410009889821040A00008",
INIT_17 => X"00401008000040300800004010000200C01000020040100802004030000002C0",
INIT_18 => X"000000C0300401008000000200C0100C01000020080000C030000000C0100802",
INIT_19 => X"325930C9A6CB261934C000200800004030040300800000020040100C03000000",
INIT_1A => X"8A28A2BD30264686668A28A2605145031C03F028000A1C2ED7831A2820244140",
INIT_1B => X"8D46A351A8D46A351AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A2",
INIT_1C => X"CFB068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D068351A",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF82B",
INIT_1E => X"54200000557FE10FFFBEAA10007FD7410FFAA97555082A800AA0000000000000",
INIT_1F => X"043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D168B55557BEAB45005",
INIT_20 => X"A8415555087BFFF55A2AA800BAFFAE9555508002AA000055574105D2A800AA00",
INIT_21 => X"087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAAA",
INIT_22 => X"0F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55A2AA955EF005568A00",
INIT_23 => X"AAA2FBD54BA080002145552ABFEAA007FC21EF007FD75FFAA8417410A2D14000",
INIT_24 => X"41000042AA10AAAABFF5508003FF55F7D568A00552EA8BEFA2AABDEAA087BEAA",
INIT_25 => X"50B800000000000000000000000000000000000000000000055042AB45F7FFD7",
INIT_26 => X"6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D5400F7A49057D08248",
INIT_27 => X"157428492E8008200043FE925571EFA380871C7028A28E3AF55F7A0925D7AADB",
INIT_28 => X"75C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA145",
INIT_29 => X"6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AAAEA8A9200249056D41",
INIT_2A => X"BE80004AAFEDB42028EBFBC2028BED152438AAA092492AAA4954281C0E2FB55B",
INIT_2B => X"FAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA007FC51C7007BD55D7",
INIT_2C => X"0041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEBAF7DF6AA00412EAABF",
INIT_2D => X"410FF84021EF0800154B20000000000000000000000000000000000000000000",
INIT_2E => X"AB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568A00FFFFEAA105D5155",
INIT_2F => X"955EF00042AAA25555410BA082E8201000043FE005D517DEBA0851574B2AAAEA",
INIT_30 => X"AAAA000804001FF005575408AA557FEB2FFAE975EF555168B55F7AA800BAF7AA",
INIT_31 => X"AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD568AA200557DE00AAA",
INIT_32 => X"07FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7D1550AAAA8002010F2",
INIT_33 => X"F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30800021EF55042AAAA0",
INIT_34 => X"000000000000000000008003FF55F7D5420BA5D2ABFEAAF7AEBDFF779A82AA43",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000200000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF0A0791B3FC1694378283C81FD996A091A32142007A336A20E03C040C002",
INIT_01 => X"A91FBDC4983088485C4A60000C24C26041280A00084000C8C212812EE2953231",
INIT_02 => X"C809AD5EB118E640A4F548FC011FF0002080000082ECC66609DB7DDDCB1FA036",
INIT_03 => X"4A120E4D3E4C90D294A31E824A52847A0B20640A88800000B8E0FD522885500E",
INIT_04 => X"001440849A2604001934800041110A71E2B068B110DB321C662AE22DC08A3448",
INIT_05 => X"370C14CA0E0800022446011C4E7F17907BEBD1AA65AE10571450DFC152522449",
INIT_06 => X"07319A109D129D450A846FE4E24C0305A1A5901C82416D05417118630839B88A",
INIT_07 => X"A5B56AD5A718C038AFFEA9FE39348C9204C389672407EE120EA5806E6C503AC5",
INIT_08 => X"C05896372728FF8C420619000003AFF4AD52A2C5D26F0EABCC96CD7AC4639902",
INIT_09 => X"5BD3571182080C000041080300F6F0C72221889C6FE20395A013282002B029F8",
INIT_0A => X"A23D203042444124098516CE0C2D13512410AD3CF8014005902DA6B2D1A4D810",
INIT_0B => X"645528937D5A85D3C4B0F883C10C24E0022B0E310612C2684CA16320A60A1185",
INIT_0C => X"288E3388E3208E3388E3288E330471904719C31438D04930ACE40FFD727C4304",
INIT_0D => X"8297A454544032252811E4AC2387F91008839C6CC413958D38C4E3208E3308E3",
INIT_0E => X"7FE0627FC25847C421516685844480204211200810028C38089AE00C894AA201",
INIT_0F => X"5D65E1E3C037E37FC3E0017C1F8037E37FC3E0017C1F900040261083080610CA",
INIT_10 => X"118796FE0037EA7FC3E0017C1F8037EA7FC3E0017C1F9300DFFFDE15D06101C5",
INIT_11 => X"BE34F00C0270F3754F1F8207FDBEBE25E0700463E17F3C7E054FF7BE6CD381C0",
INIT_12 => X"C090626DE40150459759573BBD6EF37D523E6030061341F07FC570F8FA00DFFF",
INIT_13 => X"6FE2AC3082636F301BFFFC07E00007E03F7263D383B7D1D6184131B7C1FEF64E",
INIT_14 => X"FFA0F0E06101C53E36E3D3EC84FDDDA8381C0098E57D923FDFC8D8120C4DBE0B",
INIT_15 => X"6FDF58DBF81C072540049707E0FE7323D3E43BFFF61478040570EED58F4F9397",
INIT_16 => X"00C108901822490448260224000040FC390250A2110B8ACC48B206A159A74FAB",
INIT_17 => X"08422080210882108C220842008821088230842208C20088210802308C2008C2",
INIT_18 => X"8422080230882108823080230842008C22084220842008C20080230802108C20",
INIT_19 => X"1092596D34924B2DA6884220842008821080230802108821084220842208C200",
INIT_1A => X"BEFBEFB7F7FE7EFEEE79E79EFAF2DDA73FBDCEDBFF9D3F0FDE0DB6DBF4208506",
INIT_1B => X"F77BBDDEEF77BBDDEEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"FED7BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF804",
INIT_1E => X"A800AAAAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF0000000000000",
INIT_1F => X"7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007FD7410FFAA97410082",
INIT_20 => X"A843DF55FFAA955EFA2D168B55557BEAB55005542000007FD74000055574BA5D",
INIT_21 => X"5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFFA",
INIT_22 => X"0F7D57FEBAFF80174BAAAD1555EF5555555550055574105D2A800AA00043FEBA",
INIT_23 => X"BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE95555080028A00A2FFFDE0",
INIT_24 => X"AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420BA5D2E821FFA2D5554",
INIT_25 => X"DFEF00000000000000000000000000000000000000000000000517FE10AAAAA8",
INIT_26 => X"D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC7010BEDF524AA5571F",
INIT_27 => X"1D74380851524BA5571D757DB6D5525EF555178F6D145178E00EBFBE8A101475",
INIT_28 => X"0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA147",
INIT_29 => X"92E8008200043FE925571EFA380871C7028B6AEBDF45B68A28B6DEBDF6DBEF1C",
INIT_2A => X"080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF55555057D1451524284",
INIT_2B => X"A552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45BEAA800AAFFAA9557D",
INIT_2C => X"0008517DE00AAAEA8A9200249056D4175C50920875FDA381C209256DFFDF420B",
INIT_2D => X"400F7FBC00BA55557DFF70000000000000000000000000000000000000000000",
INIT_2E => X"8A00AAFFEAA105D5155410FF84020AA0800154B2AAAA975FF5D7BC21EFF7FBD7",
INIT_2F => X"EABFF0051400A25551554BA0051400BA5551575EFF7D1401FF5D5568BE755556",
INIT_30 => X"AAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F78400145AAFFFFFEF5D7F",
INIT_31 => X"55421E75555400BA082E8201000043FE005D517DEBA0851574B2FFAABFF45FFA",
INIT_32 => X"7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF8002410FFD5575EF55",
INIT_33 => X"5D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7FFAE975EF555168B55F",
INIT_34 => X"000000000000000000000557DE00AAAAAAA000804001FF0055554088A557FEB2",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000C00000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000400322120040B313301C4389B2082",
INIT_01 => X"A74041CA38396849188160000C42424041000000090800090210090008110200",
INIT_02 => X"080108200C1000004465580000C0080100000000010432400800800009882050",
INIT_03 => X"080200010C234040842248600210812183806504488000103080014E88810000",
INIT_04 => X"0040504288A68210003120000000001002A0E8A910A072101000400A00203040",
INIT_05 => X"2800000400241801A52500094A02022014100128005004020010A1C044C02800",
INIT_06 => X"232000044084804914CA7C011AA3FC012122104CC0812D403280182308294000",
INIT_07 => X"2181020423488002940C0401D0480112000100004404004602447F8051223912",
INIT_08 => X"004812130160008304000000000021F020408264000108A00004400030400000",
INIT_09 => X"419102010104000A100348037F0584230A902A894008090343108802000FF407",
INIT_0A => X"B22D77C12052522400000400883011210000220006FC5FA400401484002447E0",
INIT_0B => X"60422291504420D084B0502044811428222300004611C57849A0150CA98A8561",
INIT_0C => X"1025B1025B0825B0825B1825B1112D8012D803003AD0413424E4014D627C0704",
INIT_0D => X"4404074040900B300A00810001A0021825E0886C0110916C96D15B0025B0025B",
INIT_0E => X"001E0800122100120499210A04A54652A12850962945180A14B44002CC020080",
INIT_0F => X"008ABA0030202100000001402068202100000001402067401026000000000031",
INIT_10 => X"00000341E8202800000001402068202800000001402062840000800000000000",
INIT_11 => X"8000000000000083D00052000100800000000000008CD0018400001200000000",
INIT_12 => X"800000069A48584000A0400000000005000000000000000048128D0002840000",
INIT_13 => X"80402000000034C1E000040000000000400FE000644000900000001A34000008",
INIT_14 => X"00003000000000004BA000112B0000880000000000807E80010010000000D1A4",
INIT_15 => X"0020250000040100000000000010CCE000198000020000000000010F80006028",
INIT_16 => X"0A728CA8C22540444924050CA9120603E0A2024048400010298432A002A00050",
INIT_17 => X"94E519465094A53946519425094A53946509425294E53946509425394E539625",
INIT_18 => X"425294E509425194E5294A519425094E5394A509465194A5294A519465094A52",
INIT_19 => X"3B1C618E38E38C31C71425294E53942519465294A53946509465394A50946519",
INIT_1A => X"8E38E39DB3B676F66EFBEFBEFAFBC5E73FC7F87A7D4ABFE7CFAFBE7BFA05004A",
INIT_1B => X"7F3F9FCFE7F3F9FCFE38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E3",
INIT_1C => X"6B23F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"00000000000000000000000000000000C0F007FFFFFFFFFFFFFFFFFFFFFFFC08",
INIT_1E => X"FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF0000000000000",
INIT_1F => X"AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFFBC0010AAD5574BA557",
INIT_20 => X"0557FE10FFFBEAA10007FD7410FFAA97400082A800AA08515555508043FE00F7",
INIT_21 => X"A2D5575EF55517FF55A2AA97400552AAAB45082E80155F7D1575EFFFAA955550",
INIT_22 => X"0FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD74000055574BA5D7FD7555",
INIT_23 => X"BAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000003DE1",
INIT_24 => X"B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE10AA803FE105D516AA",
INIT_25 => X"25FF000000000000000000000000000000000000000000000AAAEBDF45A28428",
INIT_26 => X"C7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49256DEB84104BAFFD15",
INIT_27 => X"B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE9756D145B401FFFFFF",
INIT_28 => X"DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A4904380824850381C5",
INIT_29 => X"851524BA5571D757DB6D5525EF555178F6DAAA495428412AAFB451C2A8017DE3",
INIT_2A => X"0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA2F1C50381471D74380",
INIT_2B => X"0A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D",
INIT_2C => X"00B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFFF1C7BD057D1C71FFE1",
INIT_2D => X"1FFAA84000AAFFD1401E70000000000000000000000000000000000000000000",
INIT_2E => X"75FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFDF55F78017400F78000",
INIT_2F => X"020AA0800154B2557FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2AAAA9",
INIT_30 => X"ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFFEAA105D5155410FF84",
INIT_31 => X"D5554B25551554BA0051400BA5551575EFF7D1401FF5D5568BE7AA80174AA082",
INIT_32 => X"AFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2AEA8A10082EA8BEFAA",
INIT_33 => X"557BC01EF55557DE00AA842AA0000516AABAFF8428BE7AAAEAAB55F78400145A",
INIT_34 => X"0000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000900000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0048201002842002C024500188000003000000003302300C018180006",
INIT_01 => X"020008402008404C042080000211024840000000080000080200010008110200",
INIT_02 => X"4801082248100000444008000080000041000000002222400800000009008010",
INIT_03 => X"0802010288A1484000020A400000002902006480088000003080040408810000",
INIT_04 => X"00004804890640004032030010000010008060E4100000140004500800403040",
INIT_05 => X"20000004004208016606010A0A20022000000000004000228010010080882000",
INIT_06 => X"030060004084004820906D311080020101000000008008011000000308290010",
INIT_07 => X"2100000023008002940C04000A4A010200018920646C10C50350002442003820",
INIT_08 => X"084812130160214204000000000121F000000244000100AA0004400920400000",
INIT_09 => X"419122810000081A00876882000590081100448A1000002350100CAA20002800",
INIT_0A => X"050280020100020400011640CC72602900044280028180242008069081244010",
INIT_0B => X"00200411508500B08805054C18024432A002400C99E410000080451100070014",
INIT_0C => X"05448054481544815448154481C22406A2406851201000200484950500F0145E",
INIT_0D => X"0144414A40000022880081511180036040044A013268E1205202480544805448",
INIT_0E => X"6000600010000020001102080102048102408120402800086098480008A20000",
INIT_0F => X"A2081210380021000001E003C0580021000001E003C042283426000000000021",
INIT_10 => X"00706801980028000001E003C0580028000001E003C044840000800009864038",
INIT_11 => X"80000330C00F0C0210807000010080000581C01C1C009201C000001200001607",
INIT_12 => X"8C2419101028D00020A2000000000005080082C180603A0E002A090404840000",
INIT_13 => X"8040204321188095F8000400061E001F800C202077C0009021908C4029F00008",
INIT_14 => X"00003009864038C10820201FAB000088026130071A00613E010011848322014F",
INIT_15 => X"6520350000640912058100F81C0108A0201FBA0002008239020F100880807BB8",
INIT_16 => X"114400C0002140144C2480200000040024A28400800044222980300CC4A0805C",
INIT_17 => X"2048120483204802008020082200812048120481200802008020081204812048",
INIT_18 => X"0880204812048020080200812048120080200802048320481204802008220080",
INIT_19 => X"2C208200010410400020C81200802008120C81204802008020C8120481200802",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000002A1050A",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"9840000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF818",
INIT_1E => X"5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04155550000000000000",
INIT_1F => X"AAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAAA97555F784174BAF7D",
INIT_20 => X"AAE955450055421FFFFFBC0010AAD5574BA557FFDFFF5555555EFAAFFFDFEFAA",
INIT_21 => X"A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00A",
INIT_22 => X"FA28000010552EBDE00007BEAAAAA2D14000008515555508043FE00F7AA97555",
INIT_23 => X"55557BD55FF00557FE10FFFBEAA10007FD7410FFAA97400082A800AAF7AE975F",
INIT_24 => X"B45082E80155F7D1575EFFFAA955555D51574AAAAFFD5545087FEAB455D516AB",
INIT_25 => X"7555000000000000000000000000000000000000000000000A2AA97400552AAA",
INIT_26 => X"9256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E1",
INIT_27 => X"B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7BFFF55FFA095482B6A4",
INIT_28 => X"2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF415",
INIT_29 => X"C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49003AFEFEBFBEAA001C",
INIT_2A => X"082485038F7A4905C7A28A070384120BDE100075EAA82BEDB470101C5B5057D1",
INIT_2B => X"5087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A101475D5400F7A490438",
INIT_2C => X"00AAA495428412AAFB451C2A8017DE3DF525FFFFA49756D495150492BEF1D255",
INIT_2D => X"A00555168A10002E9754D0000000000000000000000000000000000000000000",
INIT_2E => X"DF55F78017400F780001FFAA84000AAFFD1401E7FFAA97555A2AEA8A10AAD568",
INIT_2F => X"C00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215D557BF",
INIT_30 => X"028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7BC21EFF7FBD7400F7FB",
INIT_31 => X"FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2007FE8BFF080",
INIT_32 => X"D5155410FF84020AA0800154B2FF8402145A2AA954AA00043DE0000516AA10F7",
INIT_33 => X"005140000FFD140145007FE8BEF557BEAB55087FC215D555568A00AAFFEAA105",
INIT_34 => X"0000000000000000000AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"A140084000080048040100000202024040000000180800080200010048110204",
INIT_02 => X"080108020090000004655C000080000051000000002402400800000009008010",
INIT_03 => X"0002000100300C408422420002108108028065844880001030808D4288810000",
INIT_04 => X"0002584288A2C210003103001000001002A0E8C910A032541000090A00643040",
INIT_05 => X"2800080400645049A725010942220020140001A9005000004810A0C0044D2800",
INIT_06 => X"630400041404B141345A7C00426FFC01292214444081254102801A2308214004",
INIT_07 => X"21810204214080069408000008C3010200018920E06C0000021DFFA453263D32",
INIT_08 => X"084010110120018024000000000021F020408264000000080004400802400000",
INIT_09 => X"51B1004100040898128768820045142B0B902E895008080A1B13848A20002800",
INIT_0A => X"522920032052520400011641C460010D000000C8040100260008061081204010",
INIT_0B => X"4262229150012080102500211C81142880224000400411784920410C208514A4",
INIT_0C => X"0020000200002000020000200011000810008A55201000200484950004F0145E",
INIT_0D => X"40284301481509004885900101A0020964240109011890008011001020000200",
INIT_0E => X"0000200002210A320489000005A142D0A16850B6294D100A34B05242401340B4",
INIT_0F => X"00800008100001003C1FE00020080001003C1FE0002004401424008208041001",
INIT_10 => X"00000100080008003C1FE00020080008003C1FE000200080000001EA2F9EC000",
INIT_11 => X"01CB0FF3C000008000201000000081DA1F8FC0000080110080000002132C7E3F",
INIT_12 => X"3E6C00020040480040200000001004862CC19FCF81E000000010000200800000",
INIT_13 => X"004C11CF60001018000003F01FFE00004000000420800688E7B00008042000B8",
INIT_14 => X"000F251F9EC00000400004050002005D47E3F00000800084011607AD80004021",
INIT_15 => X"0000822406E5B85A3F830000000080000405000009AB87FB0000010000103000",
INIT_16 => X"1A768C68D260001448242704B912040002200640484000110104300042002018",
INIT_17 => X"B46D1B46D1B46D1B46D1B46D1B46D0B42D0B42D0B42D0B42D0B42D1B46D1B66D",
INIT_18 => X"46D1B42D0B42D0B42D0B42D1B46D1B46D1B46D1B42D0B42D0B42D0B42D0B42D0",
INIT_19 => X"200000000000000000346D1B46D1B46D0B42D0B42D0B42D0B46D1B46D1B46D1B",
INIT_1A => X"9E79E7B7F11E66C6FAD96D96520145052A1F5E2BD085122ED48F3AEB20840442",
INIT_1B => X"1F0F87C3E1F0F87C3E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"A6D4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF805",
INIT_1E => X"415555080000000087BEAA10F7803DE00FFAEBFFFF0800155FF0000000000000",
INIT_1F => X"80154105D7FC2145005155555F780155EFAAAEA8ABAAAFBFDE0055556AA005D0",
INIT_20 => X"87BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF552AA8AAA557FC0010F7",
INIT_21 => X"5D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF0",
INIT_22 => X"AAAAAA8B55F7D140010552E821EFAAAABDF555555555EFAAFFFDFEFAAAAAAB45",
INIT_23 => X"45557BE8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF5504000A",
INIT_24 => X"FFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F78402155AA8028A00A2D57FF",
INIT_25 => X"75D7000000000000000000000000000000000000000000000557BFDFFF55003D",
INIT_26 => X"FAE105D556AA10410E17555080E000280071E8A00EB8E3FE10F7AEBAFFF080A1",
INIT_27 => X"EA8AAA5571C2000FF8A17400557FC015514555757DFF8E175C7A2AAAAA82A2F1",
INIT_28 => X"FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF492",
INIT_29 => X"AF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A38492ABDE10EBDF7AF6DE3",
INIT_2A => X"5571FDFEF550E00082B6A0AFB55F7D1420104124821D7AAA0BDF6D415B575D7A",
INIT_2B => X"DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FFFFFFC7010BEDF524AA",
INIT_2C => X"00497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA001C2EA8A00F7800017",
INIT_2D => X"E00F7AEAABEF082E955450000000000000000000000000000000000000000000",
INIT_2E => X"7555A2AEA8A10AAD568A00555168A10002E9754D082E820BA08556AA00AAAABF",
INIT_2F => X"000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC21555D51575EFFFAA9",
INIT_30 => X"ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F78017400F780001FFAA84",
INIT_31 => X"843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215DA2FFE8ABA082",
INIT_32 => X"7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FFD540000000402145AA",
INIT_33 => X"5D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10AAAA975FF5D7BC21EFF",
INIT_34 => X"0000000000000000000007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000400000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000006",
INIT_01 => X"000009801830084C182060000C104268413C0A61590001D90213C10008110200",
INIT_02 => X"680108200010000054400C000080000041000000010002400800800009082011",
INIT_03 => X"0008000004002040000200100000000042800504488000103081880008C00000",
INIT_04 => X"00005042802A82100010030018000010000040C0100040140080040800003100",
INIT_05 => X"2000200400245001012100006002082000000000004000002010000040002000",
INIT_06 => X"2320400004040040144A7D000180020101000009808000000800001008210000",
INIT_07 => X"6100000021808000940800001800010200018B20206C01020200002441223C12",
INIT_08 => X"184010110120000004000000000061F000000244000081180004400000400000",
INIT_09 => X"4111002100040010008528820005100000900280000001000550860020002800",
INIT_0A => X"0080200520B23204000116404470900100402000000100242048025481024010",
INIT_0B => X"400000115040008002200000048034000002000000010712000000800F08A505",
INIT_0C => X"0000410004000041000400004100020000208201000000200404840284500016",
INIT_0D => X"00000120040000080000900201A0021924600088000000100100041000410004",
INIT_0E => X"60002000120002121C99024A00A14650A328519428651900142000000200A008",
INIT_0F => X"0000A20010200900000001400008200900000001400000001424008208041001",
INIT_10 => X"000002400820090000000140000820090000000140000A800000000000000000",
INIT_11 => X"0000000000000001500012000200800000000000000C10008400080200000000",
INIT_12 => X"0000000480004800002040000001000400000000000000004800010002800000",
INIT_13 => X"8041000000002401F80000000000000000025000274020800000001205D00808",
INIT_14 => X"004020000000000002900009AB00200800000000000012BA010100000000902E",
INIT_15 => X"652035000104000000000000001040100009BA000000000000000005400023B8",
INIT_16 => X"19028CA8D06540144C26832A1B0004000020024048400000090032A000000010",
INIT_17 => X"9425094250942509425094250942509425094250942509425094251946519465",
INIT_18 => X"4250942509425094250942519465194651946519465194651946519465194651",
INIT_19 => X"0800000000000000001465194651946519465194651946519425094250942509",
INIT_1A => X"34D34D1285B080201C92410480AB9A26667A46F345448020082E1C712A054008",
INIT_1B => X"1A0D068341A0D06834514514514514514514514514514514514514514D34D34D",
INIT_1C => X"2B60D069349A0D068341A4D268341A4D268341A0D069349A0D069349A0D06834",
INIT_1D => X"0000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF829",
INIT_1E => X"0155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA0000000000000",
INIT_1F => X"FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F7803DE00FFAEBFFFF080",
INIT_20 => X"780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555087BFDE00A2FBD7400F7",
INIT_21 => X"5D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA10F",
INIT_22 => X"A5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA557FC0010F78015410",
INIT_23 => X"45002EAAABA087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF780154A",
INIT_24 => X"E00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAABAF7D17FEBAA2AEBDF",
INIT_25 => X"8A92000000000000000000000000000000000000000000000AAFFE8A00552EBF",
INIT_26 => X"3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E",
INIT_27 => X"1FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E000280071E8A00EB8E",
INIT_28 => X"5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D556AA10410E17555087",
INIT_29 => X"571C2000FF8A17400557FC015514555757D5D71E8BEF147BFAE82A2DB555C71C",
INIT_2A => X"FFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A2AEADA38492EA8AAA5",
INIT_2B => X"2FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482B6A49256DEB84104BA",
INIT_2C => X"00A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D7000400155FFFBEDA8",
INIT_2D => X"B55FFAABDFEFF7D16AA000000000000000000000000000000000000000000000",
INIT_2E => X"20BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568BEF080402000F7AAA8",
INIT_2F => X"68A10002E9754D00517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00082E8",
INIT_30 => X"FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AEA8A10AAD568A005551",
INIT_31 => X"AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D51575EF555568BEF5D7",
INIT_32 => X"780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AAAE800AA552A97400A2",
INIT_33 => X"080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE00557BFDF55F78017400F",
INIT_34 => X"0000000000000000000A2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000800000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A14009821830284D182060000C10426840000000080000080200080000510204",
INIT_02 => X"0801080200100000046558040080000041000000002402400800000009008010",
INIT_03 => X"00020201040000D0842242024210810802006400088000003080054288C10000",
INIT_04 => X"0000400088020000003020002000001002A0E881108032100002000800203040",
INIT_05 => X"200000040000004924040108022000201000012800400010001081C040402000",
INIT_06 => X"030040040404804100006D2002A002012120004CC08125410200082308290000",
INIT_07 => X"2181020421408000940820001800010200018920206C01020200002440003C00",
INIT_08 => X"084010110120018004000000000021F020408264000000080004400800400000",
INIT_09 => X"511110010100008210010802004404230A000888400809000010042002002800",
INIT_0A => X"0000200000C04204000116404460910100082000040100240000000000004010",
INIT_0B => X"0AE22291404020902005002010000420A0200000400414684920410420200000",
INIT_0C => X"1120001200012001120011200011000090008840221000240484110000F05044",
INIT_0D => X"000803004C150100088480000980020000050001011890008011000120011200",
INIT_0E => X"000060001000020010010248040200010000800241000008009042404003E0BC",
INIT_0F => X"0080A00010202800000001402008202800000001402000000026008208041001",
INIT_10 => X"0000034008202100000001402008202100000001402002800000800000000000",
INIT_11 => X"8000000000000081400012000300000000000000008C10008400081000000000",
INIT_12 => X"8000000680001040002040000001000100000000000000004810000002800000",
INIT_13 => X"0001200000003408000004000000000040027000200020100000001A00000800",
INIT_14 => X"004010000000000042B00001000020800000000000801200000110000000D000",
INIT_15 => X"0000000001000100000000000010C030000100000200000000000105C0002000",
INIT_16 => X"03700080022100404D26A42EA01004002022000080000000018032A000A00010",
INIT_17 => X"0040100401004010040100401004010040100401004010040100400000000200",
INIT_18 => X"0000000000000000000000010040100401004010040100401004010040100401",
INIT_19 => X"0800000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"8A28A28D532A0CCC2A28A28A7AA344854A07F069CB8930AFD6A1AAA902A14148",
INIT_1B => X"6532994CA6532994CA28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A2",
INIT_1C => X"CC772B94CA6532994CA6572B95CAE532994CA6532995CAE572B94CA6532994CA",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF831",
INIT_1E => X"FEAABA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE100000000000000",
INIT_1F => X"8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA803DFFFAA843DF45FFF",
INIT_20 => X"80000000087BEAA10F7803DE00FFAEBFFFF0800155FF00042AB55FFD168B55AA",
INIT_21 => X"A2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE100",
INIT_22 => X"05555555EFF7FBC0145F78028A00A2D142155087BFDE00A2FBD7400F7FBFDFFF",
INIT_23 => X"FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555007FD741",
INIT_24 => X"EAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB55AAD168ABA002A975",
INIT_25 => X"8E00000000000000000000000000000000000000000000000557BE8BEF007FFD",
INIT_26 => X"38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E071D7AAFBEFB455D71F",
INIT_27 => X"42AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1E8B6D002090482B68E",
INIT_28 => X"D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D7000",
INIT_29 => X"2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD5410490A3DFD7F7A4821D7A2",
INIT_2A => X"410E175550071D54104951555D7EBF5C5155E3842AA00BED1421450871FFE00A",
INIT_2B => X"5BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82A2F1FAE105D556AA10",
INIT_2C => X"005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A38410E2ABD749516FB5",
INIT_2D => X"555A2FBFDF455D556AA000000000000000000000000000000000000000000000",
INIT_2E => X"8BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC01EFA2FFD7545AAAE97",
INIT_2F => X"AABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D56",
INIT_30 => X"EBFF45F78400155A2D57FE00552EA8A00082E820BA08556AA00AAAABFE00F7AE",
INIT_31 => X"D54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00FFFBD5400082",
INIT_32 => X"AD568A00555168A10002E9754D085155410085557555AAD557555A2802AA10FF",
INIT_33 => X"002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAFFAA97555A2AEA8A10A",
INIT_34 => X"0000000000000000000555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000008FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400986B830284D1820E0000C3642484000000008000008820009080A512220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"00080D4912E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"000048048002400048150300100002504230C8D9109032100020160880223000",
INIT_05 => X"220004440040080142020015001004A01200012840440000B01088C0005C2400",
INIT_06 => X"431018040014804920906C74B320020121210045408165445220082008211002",
INIT_07 => X"A5B1220421408004A56E840008B90D0200018B60A0650D450FC800644A0438A0",
INIT_08 => X"485816170760268E04000000000323F42C50826490640D28088445B0E0419003",
INIT_09 => X"41F1654100000818128728820024002B3B01AC9540080824CA13008820A02800",
INIT_0A => X"0000203600E06204000116C14474A3650048CE64E40100260048025481024810",
INIT_0B => X"08C32E915D9C208070042420180D24C8802000284007126A4D21262C20200404",
INIT_0C => X"31CA821CA831CA831CA821CA83165410E541085102000024040490A000D01056",
INIT_0D => X"812203360410110A4000840E3180021040465501011934A005101431CA821CA8",
INIT_0E => X"60006000101004A01811064B050204810240812241280D00200A08044290A088",
INIT_0F => X"482A01AAEC3602330CD2A02952DC3502330CB4A0318B41400024008208041011",
INIT_10 => X"0144C0155C3502330CD2A02952DC3602330CB4A0318B5600C587149B6D0141B0",
INIT_11 => X"083B6A51005956308D1E8202C436375908AA840AD4513437640F15245B455163",
INIT_12 => X"62F47B2872400044959BC42B1060F0D036B80B548523136C158878D8FE04E587",
INIT_13 => X"0A2699AAA3794392000D81852B0A050C224180062085134CD1719564E020C670",
INIT_14 => X"C50500D94C8121713C02B555101C90705D71009604140C0418CE0C378F0B2701",
INIT_15 => X"828E024D8C50965A40821568A06113801505010334AA73AA0666DAC20AD57400",
INIT_16 => X"123408C0822040544D248604B2100400100084008001D0113920060CDC06A27C",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"0080200802008020080200812048120481204812048120481204812048120481",
INIT_19 => X"0000000000000000002008020080200802008020080200802008020080200802",
INIT_1A => X"2082082815220A4A380000002A8313044020C0605885026853A1082100A00142",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000008208208",
INIT_1C => X"F070000000000000100800000000000000000004020000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF801",
INIT_1E => X"FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA0000000000000",
INIT_1F => X"2A801FFF7FFE8A10A28000000007FC2155F7D155545AA80001EFAAFBEAB45557",
INIT_20 => X"AFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2AEBFF45FFAEBFEAA00",
INIT_21 => X"FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEFA",
INIT_22 => X"5557FC2010002A80010A2842AAAA007BFFF4500042AB55FFD168B55AA8000010",
INIT_23 => X"EFFFD540000080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00557FF4",
INIT_24 => X"FEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021FF5D00154BAF7FBE8B",
INIT_25 => X"70AA000000000000000000000000000000000000000000000A2FFD741055003D",
INIT_26 => X"071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142ABDFC7F78E3FE28B6840",
INIT_27 => X"EBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007BC217DEBDB55555AA8E",
INIT_28 => X"AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92BEA",
INIT_29 => X"BDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA28A28BFF082ABAE10B6",
INIT_2A => X"080A175D708517DF7D497BC5028142A87000A28A2AA92007FF8F7D00042AB7DE",
INIT_2B => X"F5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00EB8E3FE10F7AEBAFFF",
INIT_2C => X"00B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E00B6DB6AA28A280001F",
INIT_2D => X"F55F7AABDEAAF784154BA0000000000000000000000000000000000000000000",
INIT_2E => X"01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBFFEF007BE8BFF5D2ABD",
INIT_2F => X"BDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BA087FC",
INIT_30 => X"AA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF080402000F7AAA8B55FFAA",
INIT_31 => X"7FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D5555FFAAA",
INIT_32 => X"AAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D2E95400A2AEA8A0000",
INIT_33 => X"FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA082E820BA08556AA00A",
INIT_34 => X"0000000000000000000FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000800000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702484000000008000008820009280A553231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"421A0A0012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"02004000890200001837830011998C31C09060DC104000102002140900003548",
INIT_05 => X"240000C400000001E404001F064000A00800000020480010A4100100001C2000",
INIT_06 => X"0300D800C1960C4400006E10B900020181840001008040057840001308212000",
INIT_07 => X"652428112180C03E8E5A2C800A3F018200418927E06686450FF8006460003A00",
INIT_08 => X"9840903525281D4F460409000000E3F08D1202C5C26A0719CC96CC7BF4629900",
INIT_09 => X"491175E10000041000C52882008600843001E09F0000002CF810200022302800",
INIT_0A => X"00002000030003040081164FC469227D2008CFE09A8180248009021091004810",
INIT_0B => X"00010C13499F01B33A00ACC0000F04F800000011800000000000433800000000",
INIT_0C => X"20CBC20CBC30CBC20CBC20CBC3065E1865E1000100000820040482B280504016",
INIT_0D => X"E7F3F01F40401C17E800C7FF3B80020000035780460124F16F06BC20CBC30CBC",
INIT_0E => X"00002200004005002001408400000000000000000000053A4096F80705FA0201",
INIT_0F => X"7B2C53F2FC16691DB587201EDDF4162B1DB527201EDDC46070241001000200F5",
INIT_10 => X"01D5CC9794162B1DB587201EDDF416691DB527201EDDD884272592D6246FC1B1",
INIT_11 => X"8E995D5A825DBA569F9FF02547068618CD3CC45B7863AE7EC00D4B122A67DF2A",
INIT_12 => X"CA5C33717461C045B5B182019473D19D7CCD856106F31A683621BDFC28800725",
INIT_13 => X"0A652CC8E3538BBA01624E51AA6C0469AC5493F5688532966471A9C5F6208C6C",
INIT_14 => X"41E1F5759001B4AA1853E6D5144AA9C914C8608D2724A4C4118D992B866E2FB1",
INIT_15 => X"825682D4A36C0B0B4B85112B2C4A05D3E6D5051893335EB0072AA85A4F9B7400",
INIT_16 => X"00800000082100544D248020000004001DC0800000010E7F70171401DE07EAD9",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0401004010040100401004000000000000000000000000000000000000000000",
INIT_19 => X"0800000000000000000040100401004010040100401004010040100401004010",
INIT_1A => X"249249120780800016A28A288028DCA30444409B054A88C5890486582A210108",
INIT_1B => X"32190C86432190C8641041041041041041041041041041041041041049249249",
INIT_1C => X"007592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2592C864",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF83E",
INIT_1E => X"0000AAAA843FE0008557DFFF0800020105D557FEAA00557DE100000000000000",
INIT_1F => X"AA8200000557DFFFF7AA80000082ABDF5508557DF45002ABDFFFF7803DE10AA8",
INIT_20 => X"07FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AAD5420000051555FFA2",
INIT_21 => X"F7FFE8A10A28000000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA0",
INIT_22 => X"05D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45FFAEBFEAA002A801FF",
INIT_23 => X"FFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA000028A1",
INIT_24 => X"BFF002ABDE00A2AABFE10082ABFFEF085542000000417555002A820AA08557DF",
INIT_25 => X"DE10000000000000000000000000000000000000000000000AAD155555A28428",
INIT_26 => X"BDFC7F78E3FE28B684070AABE803AE38145B78FD7000005010495B7AE921C517",
INIT_27 => X"547038145B505FFB6A487000005F7AFD7F7A482038002EBDF6D005B78F7D142A",
INIT_28 => X"2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00BED",
INIT_29 => X"BA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FFF1FDE821C003FE001C",
INIT_2A => X"F7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5D517DEAABEAEBFF7DE",
INIT_2B => X"5142082082005F7DFD7F7A482155BEF1E8B6D002090482B68E38FC7BE8A3DF7D",
INIT_2C => X"00B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FEF085F4703814001055",
INIT_2D => X"410007FEAA0055517DE000000000000000000000000000000000000000000000",
INIT_2E => X"FFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802AABA5D7FEAB45080015",
INIT_2F => X"FDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FEAB45F780020BA082EB",
INIT_30 => X"57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FFD7545AAAE97555A2FB",
INIT_31 => X"557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BAF7D1400BAFFD",
INIT_32 => X"7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA28428A105D7FEABEF55",
INIT_33 => X"087BD54AA550402145550000010087FFFF45F78402145F7D568BEF080402000F",
INIT_34 => X"0000000000000000000F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042604001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00020201926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"00104884880A4400403000004800027102A0E88110D83210642EA809C0203040",
INIT_05 => X"27000004004828032646000826080C201A008128044E00754010C9C192D82400",
INIT_06 => X"43000004080480492A946CE10320020121258044408125410270082308213800",
INIT_07 => X"A581424525408000AE2AA8002BC00D020003896020658FC4030000246E543AE5",
INIT_08 => X"4840101107200B80040210000002ABF02450A264002C80080004416800419000",
INIT_09 => X"4B531001000008001041080200B660E30B200C8840080A920651020002802800",
INIT_0A => X"0000203240E46204000516C04468C10100540034AC0100259001004010025010",
INIT_0B => X"04462E91440020905200A42209002420002800284002026A4D21758400000000",
INIT_0C => X"10000000000000010000000000000008000000000000002004040AA080504004",
INIT_0D => X"00000360401021280800E4000B800610C8410000A11210000000001000000000",
INIT_0E => X"6000600040D045E4195104D5854284A14250A12A512A8808289840084A020080",
INIT_0F => X"9E07A80948354B6E68982167061037496E683821670620681024000000000008",
INIT_10 => X"10B456587037496E689821670610354B6E6838216706220431961CA985D48094",
INIT_11 => X"186A91674011CE61403562274AA49CD594CF00039C7C414B6509DA22652138E5",
INIT_12 => X"3014780CC8604040424A5323845932E620295879818170304B2F5002C2043196",
INIT_13 => X"654B9104A328665603148895D44E0251142B42A3D8B2A5C8825194328A2E6A98",
INIT_14 => X"A6C6A465AA0091482382B17614F2202858EE300991415B45CD5306028F019451",
INIT_15 => X"08DC8047F17D1C7C3C02128E587D6A02B17605A130A4E8BF002258850AC5DC06",
INIT_16 => X"123508508220808048260604B2100C00022084809000D000393722A14000052E",
INIT_17 => X"284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A",
INIT_18 => X"84A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1",
INIT_19 => X"000000000000000000284A1284A1284A1284A1284A1284A1284A1284A1284A12",
INIT_1A => X"BAEBAEBFF6FEFEFEEEAAAAAAFBF7DDF77F9FBEFBFF9F3F0FDFCFBEFBF1228154",
INIT_1B => X"FD7EBF5FAFD7EBF5FAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAE",
INIT_1C => X"0077EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FA",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"57DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF0000000000000",
INIT_1F => X"7BEAB45552E80155AA802AB45AA843FE0008557DFFF0800020105D557FEAA005",
INIT_20 => X"82ABDF5508557DF45002ABDFFFF7803DE10AA80000AA087BD75EF087FFFFEF55",
INIT_21 => X"00557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAFFAE820AA5D55575550",
INIT_22 => X"FA2FBD7545FFD157555085140010F7AEAABFFAAD5420000051555FFA2AA82000",
INIT_23 => X"BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AAAEA8BF",
INIT_24 => X"EBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574BA557BE8A10A284154",
INIT_25 => X"ABD7000000000000000000000000000000000000000000000A2D155410F7FFFF",
INIT_26 => X"05010495B7AE921C517DE10A2DB50482147FFAF554971D0492E3F1C71C7BE8A2",
INIT_27 => X"1D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE803AE38145B78FD70000",
INIT_28 => X"A4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA1C7",
INIT_29 => X"45B505FFB6A487000005F7AFD7F7A482038AADF47092147FD257DFFD568A82FF",
INIT_2A => X"5D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000FFAAAFBFFBED5470381",
INIT_2B => X"24171EAA10B680124BAFFAAAFB45007BC217DEBDB55555AA8E071D7AAFBEFB45",
INIT_2C => X"00B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C20821C002AA92FFDF5748",
INIT_2D => X"010AAD157545F7AEA8B550000000000000000000000000000000000000000000",
INIT_2E => X"AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC00105D7BE8B55085142",
INIT_2F => X"BDEAAF784154BA5D5140145007BE8B55087BEAB555D04001EFF7AAA8B55F7802",
INIT_30 => X"FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007BE8BFF5D2ABDF55F7AA",
INIT_31 => X"AEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F780020BAA2FFD54105D7",
INIT_32 => X"AAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAAFBC0155085540000FF",
INIT_33 => X"5D042AA00F7FBD5410085568A10FF80020AAFFAABFF55087FC01EFA2FFD7545A",
INIT_34 => X"0000000000000000000F7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000CFFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"0002074F200904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000480488024000403000000000001002A0E881108032100002000800203040",
INIT_05 => X"200000040040080126060008020000201000012800400010001081C000402000",
INIT_06 => X"430000040004804920906C200220020121200044408125410200082308210000",
INIT_07 => X"A5A14285A15080008768A80008000D0200018B202067AF100A00002442043820",
INIT_08 => X"4850101105205380040000000000A7F42840A264920406080004400A00409002",
INIT_09 => X"411110010000080010010802000400230B000C88400808000211000002002800",
INIT_0A => X"0000203200E0620400011640446DA101004000002C0100240000000000004010",
INIT_0B => X"00422291400020900000002008002420002000004000026A4920410400000000",
INIT_0C => X"0000000000100000000000000100000000000000000000200404000000504004",
INIT_0D => X"0000022040100108080080000B80021040410000011010000000001000010000",
INIT_0E => X"0000600000000020181100400502048102408122412808082098400042020080",
INIT_0F => X"0040A100A42008000161C140000420080001C1C1400003201024000000000000",
INIT_10 => X"00022260042001000161C140000420010001C1C140001604E8084341CBA34048",
INIT_11 => X"2580E2B8802201014800C220A21829A302F1C024010C001124020C8C1A8A0396",
INIT_12 => X"0CA000048228404401004418012787124648157780120B8678C000801E04E808",
INIT_13 => X"072D04730000241000CB1325E78E0186030240000083B602398000120024ACA6",
INIT_14 => X"EF6F4163C480481506800004000CFD55196CB012481812049495C19400009001",
INIT_15 => X"800108B8FB61A0401200845594965000000400568D0CFB780055060500001001",
INIT_16 => X"123408408220000048240604B210040000008400800B0000090022A140068248",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"0481204812048120481204812048120481204812048120481204812048120481",
INIT_19 => X"0000000000000000002048120481204812048120481204812048120481204812",
INIT_1A => X"9E79E79FF3BEEEEEFE79E79EFAABCDA72E47F87BDF4EBAE7CFAFBEFB28200140",
INIT_1B => X"7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"FF83F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF83F",
INIT_1E => X"02ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA0000000000000",
INIT_1F => X"AE955455500155EF0804155EFAAD5554BA087FFFF55557BD54AAF7FBC01FFA28",
INIT_20 => X"A843FE0008557DFFF0800020105D557FEAA00557DE10A2AA801FFA28402000AA",
INIT_21 => X"552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400A",
INIT_22 => X"AA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF087FFFFEF557BEAB45",
INIT_23 => X"EF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA005568AB",
INIT_24 => X"555FFD168AAAFFAE820AA5D5557555002E80155A280000005D7FFDF4555517DF",
INIT_25 => X"0092000000000000000000000000000000000000000000000AAD1420AA087BD7",
INIT_26 => X"D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB4",
INIT_27 => X"E851FFB68402038AAAA955554900105FF0800175D7A2DB50482147FFAF554971",
INIT_28 => X"AAADB6D080A12410BE803AE38145B78FD7000005010495B7AE921C517DE10A2A",
INIT_29 => X"07FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2A0800BAE3F1C0092EB",
INIT_2A => X"B684070AA00516DABAA28402038B6803DE82F7F5D5410A2D568BC71C71D25D70",
INIT_2B => X"05D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D142ABDFC7F78E3FE28",
INIT_2C => X"00AADF47092147FD257DFFD568A82FFA4870BA555F5056D002A80155B6800001",
INIT_2D => X"145002AA8AAAAAFFC20000000000000000000000000000000000000000000000",
INIT_2E => X"00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFFF55FF84000AAAAFBC0",
INIT_2F => X"EAA0055517DE00A2AA955FFFF80020BAAAAA975450800001EF080417555A2FFC",
INIT_30 => X"0020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7FEAB45080015410007F",
INIT_31 => X"D56AB455D5140145007BE8B55087BEAB555D04001EFF7AAA8B555D557FE00A28",
INIT_32 => X"D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF803DE00FFD557400AA",
INIT_33 => X"082A80145F780020105D7BEAB45557BE8B45082EBFEBA082EBFFEF007BE8BFF5",
INIT_34 => X"0000000000000000000A2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000100000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"000440009282000001100000000000100220C8811080321000000228002A3000",
INIT_05 => X"200014C40000000100000000005C04A01000012A64400000145080C000422000",
INIT_06 => X"031042040804804100006EE4032002012120005540812540020008600831000A",
INIT_07 => X"21912244A14080008408880008000D0200018920206563000200002440003800",
INIT_08 => X"48501415032000800406180000002DF024408264000000080004400000430800",
INIT_09 => X"411100110000000010010802000400230A000880400808000450200000B02800",
INIT_0A => X"0000203000C042040001164044608101000000007C0100240000000000005810",
INIT_0B => X"0042229140002080000000200000040000200000400000684920000400000000",
INIT_0C => X"1000010000000000000000000100000800008000000000200404000010500004",
INIT_0D => X"00000260001001280000C4000300020000000000011010000000001000010000",
INIT_0E => X"400060000000000010010040040000000000000201000000000000004A000080",
INIT_0F => X"0000000000202100000000000000202100000000000004600024000000000008",
INIT_10 => X"0000000000202800000000000000202800000000000002000000800000000000",
INIT_11 => X"8000000000000000000002000100800000000000000000000400001200000000",
INIT_12 => X"80000000006000400080C0000000000D08120280000000000000000002000000",
INIT_13 => X"0040200000000010000004020010000000000000008000900000000000200008",
INIT_14 => X"0000308801400000000000040000008822110000000000040100100000000001",
INIT_15 => X"0000000004840717050000000000000000040000020000000000000000001000",
INIT_16 => X"023000000220000048240404A010040000008000000000000000020C40000008",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000200140",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"1420BAFF8000010082A954BA00003DFEF085155400F78428BEF0000000000000",
INIT_1F => X"843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD",
INIT_20 => X"AD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7AE95555A2FBE8BEFA2",
INIT_21 => X"5500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABAA",
INIT_22 => X"AA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FFA28402000AAAE95545",
INIT_23 => X"BA5D0015545AA843FE0008557DFFF0800020105D557FEAA00557DE10F7D1574A",
INIT_24 => X"0BAFFFFC20BAF7AEA8B45080417400FFFFC2145080015400AA802AA00AAAE800",
INIT_25 => X"DBFF00000000000000000000000000000000000000000000000516AA00A2AE80",
INIT_26 => X"50555412AA8ABAAADB40092E38E070280024904AA1C0438FD7005150438F78A2",
INIT_27 => X"A9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FFEDB55B6A080038E3DB",
INIT_28 => X"FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7E3A",
INIT_29 => X"68402038AAAA955554900105FF0800175D7E3FFEFBD70000124AA557FFDE10A2",
INIT_2A => X"1C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA38410038E38A2AE851FFB",
INIT_2B => X"0BE8E28A10AAA085082550A1057DBE803AE38145B78FD7000005010495B7AE92",
INIT_2C => X"001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A12410FFF1C017D14041040",
INIT_2D => X"B550855400AAF7AEBDFEF0000000000000000000000000000000000000000000",
INIT_2E => X"FF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA974AA0800020BA550028",
INIT_2F => X"57545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EFA2FBF",
INIT_30 => X"4020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7BE8B55085142010AAD1",
INIT_31 => X"002AAAAA2AA955FFFF80020BAAAAA975450800001EF080417555AAFFFDF45080",
INIT_32 => X"80015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7D17DF45007FE8AAA08",
INIT_33 => X"FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF7802AABA5D7FEAB450",
INIT_34 => X"00000000000000000005D557FE00A280020BAAAD140000A2AEBFFEF082A82010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000C00000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"0202115002BB10080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"2FE962000017102918900948514522CE09200C0D590569398ADBF8CC1E50E480",
INIT_05 => X"F05EA11E5600006B0800000038814B72A15B71D412E0AFD9C2990DA56FF0B55A",
INIT_06 => X"0640044150C025A0000000901A054F2C0A8030140BCC0460050690A95C8383D0",
INIT_07 => X"288500102F85203E8010D0AA9BC4800015001219D0550077373CAA8040006800",
INIT_08 => X"2064193920A2004B51400001414091EAA14881C0002701881B120203B7A80120",
INIT_09 => X"0409A02D965965200100104F2B00822512000000231520A024400800000ACCAA",
INIT_0A => X"0004B240028000342A00002FE00A3A1F06E649C005514AC40C082050010222D9",
INIT_0B => X"000A448C0082024AE50064B44000000000002A296AA000604838001980000000",
INIT_0C => X"044000440004400044000440004200022000200014808A02004200E540480212",
INIT_0D => X"0A80A5C8000102ED00440630004AD32400004000D58460018F6D3D8440004400",
INIT_0E => X"12AA28AA890BA00000024800480000000000000200802151025062C0BB400014",
INIT_0F => X"54E11C596A64003195933741477264003195555B418687E35836020814004049",
INIT_10 => X"99CF47DCB264003195933741597264003195555B4198843940076D296D0031F5",
INIT_11 => X"58486A556489347FE5F409CBC1362510695B6288743123C95251852041CD50A4",
INIT_12 => X"EAE2992046EB70026486035600CEC45CBCA809654B48163CCC895E1E043D4007",
INIT_13 => X"3A242DEA151848302BFD6D522B10C7EC71F6C1DB071D1216E078C4C1B1C74424",
INIT_14 => X"DAAABC982BE22267A2E2E4F44AA1DC5E37400C9EE1B7B638E8849D23C383298E",
INIT_15 => X"015998B28654565A003F0068E35352C1CAE48BFBF3A6C9B7B286B4DA8B93D037",
INIT_16 => X"009000040A8000452110A8442040D655602A102A0027E2C42320284086E6A2EE",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"1451451E96F2FC3C34F3CF3C2AC688AA263486D3260E34C0C3A7B451B0200000",
INIT_1B => X"7A7D1E9F47A7D1E9F4D14D14D14D14D14D14D14D14D14D14D14D14D145145145",
INIT_1C => X"0007D3E9F4FA7D3E8F47A3D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F4",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA0000000000000",
INIT_1F => X"80175EF0004000BA552A821FFFF8000010082A954BA00003DFEF085155400F78",
INIT_20 => X"2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D2E975EFF7D568BFFFF",
INIT_21 => X"AA8015400FF84001EF0000020AA5D00154005D043FF45555540000082EAABFFA",
INIT_22 => X"F5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555A2FBE8BEFA2843DE00",
INIT_23 => X"FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF557BEABE",
INIT_24 => X"4AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16ABFFFFAABFEAAFF84001",
INIT_25 => X"2092000000000000000000000000000000000000000000000FFFBE8BFF080017",
INIT_26 => X"38FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC",
INIT_27 => X"0925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E070280024904AA1C04",
INIT_28 => X"51420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB40092492",
INIT_29 => X"2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA410A1240055003FF6D55",
INIT_2A => X"BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC7557FC00BAE3AA9257DA",
INIT_2B => X"7F7AABAEAAF780051C70824851D7A2DB50482147FFAF554971D0492E3F1C71C7",
INIT_2C => X"00E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AABA08249756DF7D168BC",
INIT_2D => X"FFF552AAAAAA007BC00000000000000000000000000000000000000000000000",
INIT_2E => X"74AA0800020BA550028B550855400AAF7AEBDFEF08516AB55A2D16ABEFFFFBFD",
INIT_2F => X"A8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D04020AA002A955EFAAAA9",
INIT_30 => X"E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84000AAAAFBC0145002A",
INIT_31 => X"7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EF0800174BA002",
INIT_32 => X"85142010AAD157545F7AEA8B5500557DF45552A82000007BD74AAF7AEBDF455D",
INIT_33 => X"0804155FFF7D568B55FFAAAAABAFF8415545000015555A2FFC00105D7BE8B550",
INIT_34 => X"0000000000000000000AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000400000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"5295B6957FCBE0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"6DE90201BF90102103AF158E805428249851BFB2C106592088DBF8400A5055C2",
INIT_05 => X"403DA038338041EE341036BF36812841A19B68F40A807ED9C18114956FF081DB",
INIT_06 => X"00A0E2D7D3EAFF15800100FBFB333C1CBC303163670497AFF00291B3C0E20150",
INIT_07 => X"51C581123AEE54DE8008B719E61C10BBA5DAAFA9DDA1194D51E067BB00000000",
INIT_08 => X"0320A9392083056C2270E004400091181168C4D14002A110C902481FC0B42124",
INIT_09 => X"C51DFFC40C30E5F0182D0950190C0810BE00E9A76E4C6FFBE4700000B3038067",
INIT_0A => X"F7BC81C003C001674BB55B5FBB4BB4F26A19F70027CE86F047BEF19B6D94C1C1",
INIT_0B => X"0018CFC7429F326B9E822FFC00074D5A0AB033A3F330802966F74BFF8FCFB1F1",
INIT_0C => X"3EF3D3EF3D3EF3D3EF3D3EF3D3EF9E9F79E9E00185C44B91BC1740B7605040BE",
INIT_0D => X"CFEB69FF7A5F5AFFCCA787743FE67C21800367A28FC1AAF5CF6F3D3EF3D3EF3D",
INIT_0E => X"F99FD0678B87A0003000D8D02E00000000000000040025D3C21463D6BFF252D4",
INIT_0F => X"221ABD9CA854DFDD64A67D42C0F054DFDD64667D42C063E57A8F7B4594BB02C9",
INIT_10 => X"AA504801F054DFDD64A67D42C0F054DFDD64667D42C07237DFE5865F6D2BF232",
INIT_11 => X"8EAE7F5AB50D0806A9A2E0DFFF47DEDC496DA3181A0CC71440F9FBC3EFBB5AED",
INIT_12 => X"C3FC95949AEFF556EF9C75E7DCF1EB1B6E6FCDC87CB35FC94B36AECF3A33DFE5",
INIT_13 => X"AF5B6AAAE594A4C0DBFDAD94AA669809809FEFAF4157ADB55572CA527056E9C9",
INIT_14 => X"33F32ADD543430808BABAF50E1A5EB4BAEA45A250202FE0ADD39387F92B29382",
INIT_15 => X"523E865D4B1293AB6B90BF2F0E30EDEFAFD0B3FBD72E9E90D20A003FBEBF41AE",
INIT_16 => X"02F840000BCE0B6F67B3F845E017C833F6AAC02B002A2EFF22D4073DE83FB669",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9A69A6A4624C3434C0EBAEBA21B9001804F6E62029749701020B88A7CC0C0060",
INIT_1B => X"0D46A341A0D46A341A69AEBA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A6",
INIT_1C => X"00046A351A8D46A351A8D46A351A8D46A351A8D068341A0D068341A0D068341A",
INIT_1D => X"0000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA0000000000000",
INIT_1F => X"7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD17FFFF552EBFE00007",
INIT_20 => X"F8000010082A954BA00003DFEF085155400F78428BEFAAD168A000004020AA5D",
INIT_21 => X"0004000BA552A821FF5D00020BA552A82000552A821555D7FEAB55FF80175EFF",
INIT_22 => X"5AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EFF7D568BFFFF80175EF",
INIT_23 => X"55A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFFFFFDF4",
INIT_24 => X"4005D043FF45555540000082EAABFF00516AA10552E820BA007FEABEF0055555",
INIT_25 => X"AE920000000000000000000000000000000000000000000000000020AA5D0015",
INIT_26 => X"7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7",
INIT_27 => X"16AA381C0A07082497FEFB6D1451471EF007BD04920871F8FC7E3D56AB6DBEDB",
INIT_28 => X"7BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005150438F78A2DBFFBED",
INIT_29 => X"7D16ABFFE38E175EF1400000BA412E871FF550A00092492A850105D2A8015541",
INIT_2A => X"AADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5D7BFAEBA4920925EFF",
INIT_2B => X"2007FEDBD700515556DA2DF50492A2FFEDB55B6A080038E3DB50555412AA8ABA",
INIT_2C => X"000804050BA410A1240055003FF6D5551420101C2EAFBD7145B6AA2849248708",
INIT_2D => X"B550000175EFFFFBEAA000000000000000000000000000000000000000000000",
INIT_2E => X"AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFDFEFF7FBFFF55A2D16A",
INIT_2F => X"400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF5551555EF087FC200008516",
INIT_30 => X"A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800020BA550028B550855",
INIT_31 => X"7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002A955EF5D2E80010002",
INIT_32 => X"AFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FFD1575FF5504175EF5D",
INIT_33 => X"557FE8AAA000415410007BFFF450051555EFA2FBC0000A2FBFFF55FF84000AAA",
INIT_34 => X"00000000000000000000800174BA002E820105D003DFEF5D51420005D2ABFF45",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000CFFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"080BA868803F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"42016B0C401F58495C900A4859552A611D9A640F5903B2388004004C08A06008",
INIT_05 => X"7008000E0E508C01C28640000801133060E0032801E0202000991B708280B501",
INIT_06 => X"560000000022229A60B048048120FF040000000002C44D620F0228454C838100",
INIT_07 => X"58800A001D4033A004904087F9E3901218050018024110D6771C1F90C2856828",
INIT_08 => X"3020A82929A807B3731021400058C020000A9729400D10100420480202AC2140",
INIT_09 => X"0419002D86184A01018030430700802541420440022030041A814A0080064C1F",
INIT_0A => X"0000F0CA8428642430080438408A510185A200000045C18C0E0000A0820500B9",
INIT_0B => X"311324AA2373088479105D044A1022000001835C0C30C2E21480349D00100202",
INIT_0C => X"000C2000C2000C2000C2000C2000610006100100180A8062026000DC425C0301",
INIT_0D => X"10108003C00021002046088B5001FB3650D89844703657083080C2800C2000C2",
INIT_0E => X"007E281F840C00284A17210001060D8306C18360C1380A0260CB980840080810",
INIT_0F => X"9BBEF8E50B041029075982BF3873041029079982BF39748AA0AC800014804032",
INIT_10 => X"79BFD7F7F3041029075982BF3E73041029079982BF3F632C5F96D3C11555D5D7",
INIT_11 => X"A595405FC7F1CFEBC7586C4100A53162B47FD7E39FFEECE1598702345156AEA4",
INIT_12 => X"FE037ACFB88083A99E06271BB0CA207DFDD5920057E0B001B0EBCC79932C5F96",
INIT_13 => X"2A002DD51B6F7FC4A411D1E8D44517F14EAFE36E55150016EA8DB73E39464006",
INIT_14 => X"C30351452A13D55CFFA76E928E3891F148B30399F5FB7F28C800DFA06F5DF5CA",
INIT_15 => X"57DFEAEF1005475F1D1F608819CF0EE76E12C824ADD9089715F25FAF9DB84953",
INIT_16 => X"34041A41A0000010180C02801680460FC900052FA10DC0006DA4881C110155AC",
INIT_17 => X"60D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8",
INIT_18 => X"0D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D83",
INIT_19 => X"00000000000000000020D8360D8360D8360D8360D8360D8360D8360D8360D836",
INIT_1A => X"8A28A2891182C8A82E0820825945DF675C0770B9E11807E54587BEF8B0000000",
INIT_1B => X"2552A954AA5128944AAAA28A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A2",
INIT_1C => X"000128944A25128944A25128944A25128944A25128944A25128944A25128944A",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E954000000000000000",
INIT_1F => X"D568B55080028B55002E82000087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD",
INIT_20 => X"87FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA087FFFFFFFFFBFDF45AA",
INIT_21 => X"0051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE000",
INIT_22 => X"00804154BA55042ABEF5D7FD75FFAAD540145AAD168A000004020AA5D7BE8B45",
INIT_23 => X"10557FD7545FF8000010082A954BA00003DFEF085155400F78428BEFAA800000",
INIT_24 => X"000552A821555D7FEAB55FF80175EF5D00020105D2A97400082E95555085168A",
INIT_25 => X"24280000000000000000000000000000000000000000000005D00020BA552A82",
INIT_26 => X"E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A9",
INIT_27 => X"FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147FFFFFFFFFBFDFC7EBF5",
INIT_28 => X"003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092087",
INIT_29 => X"C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AADF6DB7DE3F5FAFC708",
INIT_2A => X"F78A2DBFFA28407038140410492550A2ABC7497BD25FFAADF4516DBED16AA381",
INIT_2B => X"8002E9557D1C516FA28417BD5545E38E070280024904AA1C0438FD7005150438",
INIT_2C => X"00550A00092492A850105D2A80155417BEFB6DEB8E175FF5D0E0500049209742",
INIT_2D => X"FEF552E974AA082A820AA0000000000000000000000000000000000000000000",
INIT_2E => X"DFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFFFFFFFFFFDFEFF7FBFF",
INIT_2F => X"AAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AA557FF",
INIT_30 => X"FFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D16ABEFFFFBFDFFF552A",
INIT_31 => X"FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087FC2000FFD56AB45A2F",
INIT_32 => X"50028B550855400AAF7AEBDFEFA280154BA550400000552AA8B45087FC01EFA2",
INIT_33 => X"5D2E974000804154BA082A975EF5D517DEAA007BD5545AAAA974AA0800020BA5",
INIT_34 => X"00000000000000000005D2E80010002A954005D2A82155087FFFFEFAAAA975EF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000400000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000010228001000000000000000000024001620280000000000354200004008",
INIT_04 => X"00016200001310090090004840004152C7208802590000388000004C08006000",
INIT_05 => X"7008000E0200000000000000000100302000000000E02000009900000000B100",
INIT_06 => X"00000000000000100000000000001B040000000002C42010010200004C838100",
INIT_07 => X"E0050A040041593104004500480090080A011202201400204204018000000000",
INIT_08 => X"30E409080188000021A0000100004082A140102B4020109801A4CE0037100100",
INIT_09 => X"00000005861840000000004301000B000000000001C1C0000000000000020C01",
INIT_0A => X"0000B0C0000000101400040C0408100000000000004540800000000000000099",
INIT_0B => X"000010000800011000000000000000000000BC0007C00008092C800080000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"08000EC0000000000000000010004B2000000000000000000000000000000000",
INIT_0E => X"0006280180040000000000000000000000000000000000000000000000000001",
INIT_0F => X"4451B81A70AB3006BA0011400760AB3006BA0011400680F02096834820000000",
INIT_10 => X"04082248A0AB3006BA0011400160AB3006BA0011400084C780687DBA82800808",
INIT_11 => X"796E80A00802301BC0A7531EDD98E73B02800804620D030F873EB49F30B80112",
INIT_12 => X"0000002044F091A860700FF9198AA115D5DA37F7A80C8A3604001C0664C78068",
INIT_13 => X"51AC9000000000314E01F9F30198600631448410A2A8D64800000081B0A936B0",
INIT_14 => X"0303842281C80A23004411AD661891F15148A4420804241526D6000000000985",
INIT_15 => X"35F3D282000C6C5456C84850F61050C411AD6284FDA861682805A04A1046B2E0",
INIT_16 => X"00000000000000000000000000004600C0013800003088004202304366A4A9D3",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"86186186851046260A9A69A6039045DD1F863808633005010063A20C90000000",
INIT_1B => X"930984C26130984C261861861869A61861861861869A61861861861861861861",
INIT_1C => X"0000984C26130984C26130984C26130984C26130984C26130984C26130984D26",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BA0000000000000",
INIT_1F => X"FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082",
INIT_20 => X"87FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7FFFFFFFFFFFFFFFFF7",
INIT_21 => X"080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA0",
INIT_22 => X"FF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFFFFFBFDF45AAD568B55",
INIT_23 => X"00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AAF7FFFFFF",
INIT_24 => X"B55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB55A2FFFDFEF5D2EBFE",
INIT_25 => X"04AA000000000000000000000000000000000000000000000AAFFFDF45A2D16A",
INIT_26 => X"FDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA00001",
INIT_27 => X"FFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7FFFFFFFFFFFFFFFF7FB",
INIT_28 => X"00001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92EBF",
INIT_29 => X"3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7F1F8FD7AAD16AB4500",
INIT_2A => X"087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D000000010087FFDFC7E",
INIT_2B => X"DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6DBEDB7FFEF552AB8E38",
INIT_2C => X"00B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E284971F8FC7AAD56DB6",
INIT_2D => X"FEF552E954AA0004000AA0000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFFFFFFFFFFFFFFFFFFFD",
INIT_2F => X"175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00557FF",
INIT_30 => X"56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FBFFF55A2D16AB550000",
INIT_31 => X"0402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AAF7FBFDFEFF7D",
INIT_32 => X"FFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7FFFFFFF552AA8BEF08",
INIT_33 => X"08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA0008516AB55A2D16ABEFF",
INIT_34 => X"0000000000000000000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000800000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"0001E6000053300B00D0005800000000000000407B0004BB830004DC3D01E000",
INIT_05 => X"F0FF433EFE022001C81080001101F977E0201C409BE1F10623BB000A100CF300",
INIT_06 => X"0F00100002E22EB440012C809B2FFF7C8E8840155FDC0000010E40087D8787A1",
INIT_07 => X"3B800000000000000008407FC800B0000000100600040000C205FF91C000F800",
INIT_08 => X"28C0B0300020852000002101554021F000000000000000090492260200002000",
INIT_09 => X"00000007BEFBC010002008FF7F00000000010018A81000041C401000004FFDFF",
INIT_0A => X"0002B7C0000008000000200000200A0C004408C2007D5FC800000240001227FB",
INIT_0B => X"000000000000000000000000800800A400000000000000008000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000800080000000",
INIT_0D => X"001000000100000020000800101FFB6000000000000000000000000000000000",
INIT_0E => X"07FE29FF800C00000001002040000000000000020480002E42429C0000080000",
INIT_0F => X"4D4E180010040000400000001E60040000400000001E6010003C000000000030",
INIT_10 => X"000094B1E0040000400000001E60040000400000001E60804000000400000000",
INIT_11 => X"02000000000033628000100100000004000000006170C0008001000004000000",
INIT_12 => X"000000295810000000A100020614148002000000000004307CC3CC0000804000",
INIT_13 => X"2000000000014AC000120200000000003F0D800020100000000000A4B0020000",
INIT_14 => X"0C0C00000000002E2D000001006204040000000005786C004000000000052580",
INIT_15 => X"0A0C0939BEE1810080200000E0CE0EC000010020000000000000AE8A00002002",
INIT_16 => X"8040400400C08080000000000049F6FFC0100000000000008008008000400010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000200",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C30C320624C1090D0F3CF3CD038001801C10000804482A60D09008269020010",
INIT_1B => X"86432190C86432190CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C3",
INIT_1C => X"000432190C86432190C86432190C86432190C86432190C86432190C86432190C",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"4174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804020100000000000000",
INIT_1F => X"FFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA000",
INIT_20 => X"87FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFFFFF",
INIT_21 => X"552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA0",
INIT_22 => X"FFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFFFFFFFFFFFF7FBFDFFF",
INIT_23 => X"EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA007FFFFF",
INIT_24 => X"FEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDFEFF7D56AB450000021",
INIT_25 => X"5000000000000000000000000000000000000000000000000F7FFFFFFFFFFFFD",
INIT_26 => X"FFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA08000",
INIT_27 => X"FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428087",
INIT_29 => X"FFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFFFFFFFEFF7FBFFFFF55",
INIT_2A => X"B6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AABEDF6FABAEBFFFFFFFF",
INIT_2B => X"7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7EBF5E8B550000071EF",
INIT_2C => X"00FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AAA497FFFFFFF7FBF8FC",
INIT_2D => X"FFF5D2A954AA0800174100000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410A2FFF",
INIT_30 => X"BFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFFFDFEFF7FBFFFEF552E",
INIT_31 => X"FFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00AAFFFFFFFFFF",
INIT_32 => X"2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAAD16AB450804174AAFF",
INIT_33 => X"087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA557FFDFEFF7FBFFF55A",
INIT_34 => X"0000000000000000000F7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"1094EC681244819000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"0001E6000053300F01D4587800446194F49020107F0012BBC00202DC3823EA82",
INIT_05 => X"F0F807BFFE000120080002341881F3FFF012412A9FE1E01013BF09404050F300",
INIT_06 => X"08808210996035A000006EC2E04FFFFC0A0000101FFE4036450E08247F878703",
INIT_07 => X"003400812A156C002822987FC830F40134CC74D002016612DE87FFE004008040",
INIT_08 => X"02348D2D00080C0C53400044114000000D022640B42406808790055043A82824",
INIT_09 => X"080AC707FEFBC110008420F7FF388B70A20389346FE8000580200800008FDFFF",
INIT_0A => X"4636FFC00080013029811240444A82422A828C03BC7D7FC15025B1AB6E85A7FF",
INIT_0B => X"2019480E63180855A492712CC01C49C20201BFE45FF0C004041DA2218A8A3151",
INIT_0C => X"648A3648A3648A3648A3648A366451B2451B210018C241102068006C620C0388",
INIT_0D => X"80050094104431200090080C621FFBE0008A94641165448C80C103648A3648A3",
INIT_0E => X"9FFEADFF8050250010030165290008800440022201082401A002000C48000201",
INIT_0F => X"48A004A6C0D2820302C005A83480D1820302A009B02B101390C0CB2830816202",
INIT_10 => X"8904831400D1820302C005A83480D2820302A009B02B021A85C0941150013180",
INIT_11 => X"8834600024D052C1051E0B92D400360520202682C19024B6164E300448510140",
INIT_12 => X"4093E22A2012418A9D1D44ADD9E0F174103820101C0B8160D5516259FA1A85C0",
INIT_13 => X"8AA288209E615100280DA0052000C5006402000206C55144104D510CC1B0D640",
INIT_14 => X"D50020C04023033C52009144231D902818100C90058010361AC808126C88660D",
INIT_15 => X"2386454988140600C0181500A13E830011008B0374007000B4E0CD00024500A0",
INIT_16 => X"0224004002000000703804008001F7FFF01B982B01258088C008CC41198A1220",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"0000000000000000002008020080200802008020080200802008020080200802",
INIT_1A => X"BEFBEFBFF7FEFEFFFE79E79FFFF7CFF77FBFFEFBFF9F7E0FDF9EFEFBF0000000",
INIT_1B => X"FF7FBFDFEFF7FBFDFEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000100000000000000",
INIT_1F => X"FFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080",
INIT_20 => X"7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAF",
INIT_22 => X"FFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFFFFFFFFFFFFFFFFFFEF",
INIT_23 => X"AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFF",
INIT_24 => X"FFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFFFFFFFBFDFEF5D2A954",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA00000",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAF7F",
INIT_29 => X"FFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFFFFFFFFFFFFFFDFEF55",
INIT_2A => X"082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA002A95400087FFFFFFF",
INIT_2B => X"FF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA",
INIT_2C => X"00E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50BA557FFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0000020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAFFFFF",
INIT_30 => X"FFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E",
INIT_31 => X"2E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410087FFFFFFFFF",
INIT_32 => X"7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7FBFFFFF552E954BA00",
INIT_33 => X"5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA557FFFFFFFFFFFDFEFF",
INIT_34 => X"0000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"8632CA211E4491D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"24B000808800040439245B221373581F97B0A8D1040F92000F42000047A00E58",
INIT_05 => X"0107C4410008816B105036B4180C000811E9BF2844021B1004045E4249500449",
INIT_06 => X"0111C2D50A46AE45281502E4A2200081ADA0E054402365774611E047020008E0",
INIT_07 => X"80BD5AA4BF5C91F840C1710010344DB9A808FDFF3DE0313014A2007540401804",
INIT_08 => X"EA212D6D481ADF0CE47CA21544009007A64EBD64049D028B93D9561A48F60276",
INIT_09 => X"0E48D500400015805060040080A2A0F4A82381B4000A0905A0283800AA500200",
INIT_0A => X"4E700838460402635019FBFE7FCA13520F8AAD050402204090090319A5002004",
INIT_0B => X"040F4A944B1AA313C0022AA0011C0DC0002800134000000849BCC3240A8A7151",
INIT_0C => X"70AA070AA070AA070AA070AA072550385503800500001840000C80B410014088",
INIT_0D => X"0A9CA0D458D131652A154CAC6B600085080B14004D1594832824A070AA070AA0",
INIT_0E => X"C00044000A1EC1C44140D101A54280A14050A028500A84F02842A24C594A0687",
INIT_0F => X"59E0C4E6C256690581800F1C3E82562B0581200F1C3F08145602280402080448",
INIT_10 => X"AB8581B602562B0581800F1C3E8256690581200F1C3F1238473F121000613383",
INIT_11 => X"0E1050083750B3E4275F829547008600C030374361FA2CEE046D48122C438100",
INIT_12 => X"C012A66F61154C019511628756231018500C00203E138061565160782238473F",
INIT_13 => X"AA612C0096C37B00D1724801A0009C606D1221D104553096004B61BCC1128C4C",
INIT_14 => X"41E0F0600035842E7601C2C4AC68A98810080AA825A890225189980254CDE608",
INIT_15 => X"637E00D0A1080301401C390320188321C2C0B13890105800D520AF94870B012A",
INIT_16 => X"22F110111B281A54753AA004002601001918008C10912A4440B24E8B58234A89",
INIT_17 => X"0882208822088220882208822088220882208822088220882208822088220882",
INIT_18 => X"8020080200802008020080200802008020080200802208822088220882208822",
INIT_19 => X"8000000001FFFFFFFFC802008020080200802008020080200802008020080200",
INIT_1A => X"9E79E7BFF3FEFEBEEEFBEFBEFBEFDFEF7F47F8FBEF5EB7E6CFEFBEFBE8289144",
INIT_1B => X"7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"0003F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000000000000000000",
INIT_1F => X"FFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFF",
INIT_24 => X"FFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFFFFFFFFFFFFF552A974",
INIT_25 => X"0010000000000000000000000000000000000000000000000007FFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0804154BAF7FFFFFFFF",
INIT_2B => X"FFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA",
INIT_2C => X"00007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000AAA2FFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804000100000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A",
INIT_31 => X"04174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAF7FFFFFFFFFF",
INIT_32 => X"FFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E974AA08",
INIT_33 => X"AAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA2FFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"5886C0201A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"0005EE040057700F40D08078500000D9218020407F0000BB8018A2FC380BEAC2",
INIT_05 => X"F0F817FFFE400800020224000405F7FFE0124002FFE1E0C517FF09111212F300",
INIT_06 => X"400000409120338860900482404FFFFC000000001FFC0832050E00047F97870B",
INIT_07 => X"00246801C41C3E81E872C8FFE900FC31348EFDF03BE15E22DA07FF92C2041020",
INIT_08 => X"6220280D2B025988311AB14155421006891A1089F6E200000022C140068EB902",
INIT_09 => X"0002021FFEFBC80000000077FF184B03010004002FE1F2900201000000FFDFFF",
INIT_0A => X"0006FFEA002020626995FBE077430001E7320006F87D7FA84024B0225A890FFF",
INIT_0B => X"241C482B20400CC52492710CC80060020A81BFE41FF0C2060481200180000000",
INIT_0C => X"040430404304043040430404304021820218210018C24110A860006C620C0312",
INIT_0D => X"001002001804800000952800001FFBF040C088669070510C90C1430404304043",
INIT_0E => X"1FFEAFFF805025E00853B92588000400020001000020A8018008002000014030",
INIT_0F => X"148484054395E27E428002A4200397E07E422002A420100382FCC30832A16382",
INIT_10 => X"788417000397E07E428002A4200395E27E422002A420110A51C01C0590401486",
INIT_11 => X"1A2490040590C08120558C1759BE1C05A0400383808800DA1929F728641100C0",
INIT_12 => X"00136006000215EA0A4833A32C8832050028603050014031B3950000C90A51C0",
INIT_13 => X"658280009A2030108B14AC05C00112405222088B8332C140004D101800CE7200",
INIT_14 => X"B6808060201281004228996085F10020180C030880D11019CE4000026C00C006",
INIT_15 => X"49DC7143F01C04240030720641E0A028996483A17204680410A04104A2659196",
INIT_16 => X"1000080080000000000002001201F7FFC0011C2F81A48080CA32800A0108152A",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"0000000000000000000040100401004010040100401004010040100401004010",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080002010FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA08",
INIT_33 => X"F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"0000745C200801000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"0001E6000053300F00D0007810042140C00000407F0000BB800000DC3801EA00",
INIT_05 => X"F0F8033FFE000000000000000001F17FE01240009BE1E00003BF00000000F300",
INIT_06 => X"000000009120110020100002404FFFFC000000001FFC0000010E00007F878701",
INIT_07 => X"00102050840950002802C87FC800FCAA035400001B918600C207FF8000000000",
INIT_08 => X"6234AD280B02500063AC2840001610020408178B600C24000136496087300042",
INIT_09 => X"00000007FEFBC00000000077FF000B00000000002FE0000000000000000FDFFF",
INIT_0A => X"0006FFE80000015406A800003388000025000002387D7F804024B0224A8107FF",
INIT_0B => X"20502000200000400490510CC00040020201BF441FF0C0000000000180000000",
INIT_0C => X"040030400304003040030400304001820018210018C0411020600048620C0300",
INIT_0D => X"800B00000000000000000000001FFBE0008080641060400C00C0030400304003",
INIT_0E => X"1FFEADFF80002080000000208800000000000000000020018000000000000004",
INIT_0F => X"009181008024A00043601100210024A00043C0110020901382CCCB28B0806202",
INIT_10 => X"040A03080024A00043601100210024A00043C01100209240C840C201D0210840",
INIT_11 => X"A604E0080820009908008341B000A8212070082002890010068320860C920180",
INIT_12 => X"00800082041205EC00044C1ACB66C37542082030281E0580001012811A40C840",
INIT_13 => X"27A004300004103160DB3005E000618040C022000593D002180002090166B406",
INIT_14 => X"FF20406040084210C062000C2A2DDD00180C04504086002CD680C0100010480B",
INIT_15 => X"04295C98F80400008040CC0582169022000C2876C404780028500160880012BB",
INIT_16 => X"0000000000000000000000000001F7FFC001B823018F00880008805241060208",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9EF9EFB263CC3090CABAEBAFF96857757B73E6089966B9EF9D5A220CC8000000",
INIT_1B => X"0F0783C1E0F0783C1EFBEFBEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF",
INIT_1C => X"0000783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2010000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020100000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA00",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00004000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"4909E6093253306F82D0007C80000000080E01007F8020BBC00040DC3801EA00",
INIT_05 => X"F0F8033FFF0240012C1400080291F17FF01241009BE1E00203BF80800000F392",
INIT_06 => X"0DC00CC0992033A062116E82404FFFFC0E0801101FFC0000010E08A07FC78701",
INIT_07 => X"00000000000000002802C87FC800F8000000000019810600C207FFF3C410D841",
INIT_08 => X"E8002000080281000008A0000014100200081000000000080480AE0000002000",
INIT_09 => X"80040007FEFBE031018C31F7FFBAEBC0020008086FE0000100280800000FDFFF",
INIT_0A => X"0006FFF800C04000000000003300800005000032387D7FE94FBEF2B2CB8DA7FF",
INIT_0B => X"20100000200000400490D10EC00040220201BF441FF0C0600000000180000000",
INIT_0C => X"04003040030400304003040030400182001821001DCCC31222730A49620C0300",
INIT_0D => X"000000000000000000012800001FFBE0008080641062400C00C0030400304003",
INIT_0E => X"1FFEADFF805025C0304001E58906088304418222C108A009A090400000000000",
INIT_0F => X"00100100000480000200100000000480000200100000100380F0C30830A06302",
INIT_10 => X"0008000000048000020010000000048000020010000000004040000010000000",
INIT_11 => X"0004000000000008080000011000000020000000020000000001200000100000",
INIT_12 => X"000000800002018C010000020800000800122000000004004000008000004040",
INIT_13 => X"2080000000040000001020020000000000800200001040000000020000021000",
INIT_14 => X"1000008001000000800200000021000020100000000200004200000000100000",
INIT_15 => X"0008400000000605000000000200000200000020400000000000002008000002",
INIT_16 => X"226410410346010000000400A011F7FFE0031823010400800000800001840000",
INIT_17 => X"2088220882208822088220882208822088220882208822088220882208822288",
INIT_18 => X"0882208822088220882208822088220882208822088220882208822088220882",
INIT_19 => X"17FFFFFFFFFFFFFFFFE088220882208822088220882208822088220882208822",
INIT_1A => X"0492410A048029890AD34D35FDD144A50CB5462D14997BE09E760AED04040000",
INIT_1B => X"6231188C46231188C49249249249249249249249241041041041041041049241",
INIT_1C => X"000B158AC562B158AC562B158AC562B158AC562B158AC562B158AC562B1588C4",
INIT_1D => X"0000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"94A7B2B1450000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"6FEBEF5FEC737AFBC6F85FDEB220109E1FEFFFE3FBA7FDFB9BD301DC3FF5F0D2",
INIT_05 => X"F0FFEB3EFFF7FDED3FBFF6A84383F177F5FB7FF59BE1FF980BBBB7FE6D21F3DB",
INIT_06 => X"FBE564C71268F3BBF5FBFC2A427FFF7C3E3A74667FDDB7FB870FF30FFDEF87F5",
INIT_07 => X"3BC18306396FBEC14489737FDC00B13BB79DFDB83BF4112AF205FFBDD3AFB93A",
INIT_08 => X"21E4391909B381B0B1F8E041051831FA3068D77E000030021324620C0B9C2060",
INIT_09 => X"D13D980FBEFBEBF30B8D79FF7F451F33CFD60FE8FFFDF54003B1D4223B4FFDFF",
INIT_0A => X"B5AFF7CFACFAFE776F39FF7077E29D83CFAB300B017F5FFE6FBEF73BEFB967FB",
INIT_0B => X"737AF3FD62601EDC25B3533DCEB07F262213FFC67FF1C7FBFB5EC9478D5DA3A3",
INIT_0C => X"5E3035E3035E3035E3035E3035E981AF181AE315BDDCC3B336F7C548667D47B7",
INIT_0D => X"100C0E60FB9FC3A80EF69A004DFFFF7FF5F9A06E19F4DA0E80E903DE3035E303",
INIT_0E => X"7FFFF9FF8FAFAA3ADEBFB9726BAF5FD7AFEBD7F7EFFD7ACDB7F947F0EA035CF6",
INIT_0F => X"0080A40403E8BD8002000FC02003E8BD8002000FC02010979AFFE36C36B86702",
INIT_10 => X"EE00034003E8BD8002000FC02003E8BD8002000FC020037B0040A00010003E02",
INIT_11 => X"C00400003D80008160400FD81341C00020003B80008C00801EF0285380100000",
INIT_12 => X"81038406809677FA080468C46A81080581002000780C8001C8100201037B0040",
INIT_13 => X"90D162001C803411FC0024080001F80040026C0807C868B1000E401A01F11909",
INIT_14 => X"10503A00003E020042AC080CEB01228A80000F600080123E232130407080D00F",
INIT_15 => X"7520750001064180807868000110C02C080CFA0042400000F8800105B02013F8",
INIT_16 => X"FF7EFEEFF3EEC3FF7FBFFBCB7FFFFEFFE00BFF7FEBF420800EC0CBEE61F81008",
INIT_17 => X"F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F7FD",
INIT_18 => X"5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7",
INIT_19 => X"37FFFFFFFFFFFFFFFFF5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F",
INIT_1A => X"A61861BAF15EAA6AFC38E38EA3AD8ADE7A48F0B366429F434AA9FC376DAE4432",
INIT_1B => X"130984C26130984C261861861861861861861861861861861861861861869A69",
INIT_1C => X"0000984C26130984C26130984C26130984C26130984C26130984C26130984C26",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"1085B0B041000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"6FAB975B6470BAF386C87A9CB00000001FEF9F23E3A7BDE79B5101D23FB5C0C2",
INIT_05 => X"C8FFCB38FF35B44C25ADE72041A3F147F5FB7F759B91FB880BA3B6FE2921CBDB",
INIT_06 => X"B98420C71408D113956AFD0842FFFC7C3032646EFF1DB7FA868FE30EF1CE47E5",
INIT_07 => X"0041830600640C415004637FC4003021259CFDB01BF80028E001FF8251AB9D1A",
INIT_08 => X"200822020842203000082050000110023068D030000028200000008400000051",
INIT_09 => X"90A4880E3DF7E2FB0B8E717C7F411F3BC6D60B60FFDDE440018AC4AA3B0FD1FF",
INIT_0A => X"042787C5AC5ADC424B39FB6073D00D8048A31008017C1F826FFEF41FEEB027E3",
INIT_0B => X"7BEAF1C152201A4C05B7531D56B05B06A213FF863FF5D5F9FB5E8847A0702606",
INIT_0C => X"0D1030D1030D1030D1030D1030F0818688186B51BFDCC39732F3554866AD57C3",
INIT_0D => X"10080A20ED1D41880CC61A0044DFFC6EB5BCA06F18FC5A0E00F0038D1030D103",
INIT_0E => X"3FFE91FF98AEAA1AC6AC9A3A4AAD5B56ADAB56D5AFD572C597B147506203E8FC",
INIT_0F => X"0000260403C8948002000EC0000BC8948002000EC00010878AC3CB8AB8857202",
INIT_10 => X"EE0000400BC8948002000EC0000BC8948002000EC000097B0040200010003E02",
INIT_11 => X"400400003D80000070400DD81041400020003B80000410801AF0204180100000",
INIT_12 => X"010384008086378A080428C46A80080081002000780C800188000301017B0040",
INIT_13 => X"909042001C800409FC0020080001F80000007C0807484821000E400205D11101",
INIT_14 => X"10100A00003E020000BC0808EB01020280000F60000002BA222020407080102E",
INIT_15 => X"7520750000024080807868000100403C0808FA0040400000F8800001F02003F8",
INIT_16 => X"EF3AF6AF6389C2FE128971AB2DDDF8FFE0031B776BF4208006C0C92621F81000",
INIT_17 => X"D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B5",
INIT_18 => X"5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56",
INIT_19 => X"3FFFFFFFFFFFFFFFFFD5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D",
INIT_1A => X"0000001E0080397908000000A48710B4080240E543021B438A010825238B443A",
INIT_1B => X"4020100804020100800000000000000000000000000000000000000008200000",
INIT_1C => X"000A05028140A05028140A05028140A05028140A05028140A05028140A050080",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"8C2100804900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"02000100440408002408008002221000204116A280000F000001400000100010",
INIT_05 => X"00000000001265050080C000190002000000005C0000000A0000002C20600000",
INIT_06 => X"14016012000C405280200008001000011110012220009A88800009A880000000",
INIT_07 => X"0048912242288100800102000400010208000000040000082000002400814008",
INIT_08 => X"0A010040401080308400821155540001122448142491008A0049120408402210",
INIT_09 => X"04080A000000124058200408000880004440004080160C4100A8580099400000",
INIT_0A => X"4A50000080080E041000000008000C81000110010500002000000180001C8000",
INIT_0B => X"110091500020B408810000100200020408B0000020000081B2C208420ADA5353",
INIT_0C => X"5814058140581405814058140580A02C0A02C004800210C19808400500010009",
INIT_0D => X"10040860B188C0A80653020005A004039010280000800B00100040D814058140",
INIT_0E => X"600010000280000802050010660001000080004004900204020105302A000C42",
INIT_0F => X"0000A00000081480000001400000081480000001400000800C01082082210500",
INIT_10 => X"0000024000081480000001400000081480000001400000010000200000000000",
INIT_11 => X"4000000000000001400000080041400000000000000C00000010004180000000",
INIT_12 => X"0100000480802A40000000400000080081000000000000004800000000010000",
INIT_13 => X"1010420000002400040000080000000000024400000808210000001200010101",
INIT_14 => X"00100A0000000000028400004000020280000000000012002020204000009000",
INIT_15 => X"1000000000024080000000000010400400004000004000000000000510000040",
INIT_16 => X"8408420430E699AA42A1508104EA08000000810020000000044001AC20500000",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_19 => X"8000000000000000000010040100401004010040100401004010040100401004",
INIT_1A => X"20820800D41A8283AC618618EF1088160885001234B96061CCDEC4D205061170",
INIT_1B => X"6030180C06030180C08208208208208208208208208208208208208208208208",
INIT_1C => X"000B0582C160B0582C160B0582C160B0582C160B0582C160B0582C160B0580C0",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0803B2814D0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"26E1E905CC574828C4F85FC600000016004F77E2F887CDB80BC340DC07D1F000",
INIT_05 => X"F007E33E01D26CE43A92F2880B01F37011E93ED49BE01F1A03B8972E6D20F049",
INIT_06 => X"5AA06002026872BAE0B1282A005FFF001E1870223FC3BFC98101F109FC6780F1",
INIT_07 => X"3BC081023B233E804488527FDC008019968D74982C94110AF204001BC285A828",
INIT_08 => X"01E4191901A101B031F84000000831FA1028575A000110800124600C039C0020",
INIT_09 => X"C1111A0782082B50080508FF00048B124D4005C8AFF4154102914800110FFC00",
INIT_0A => X"B5AAF00A80A82C332D18ED301D229C82C7A93002017F405C409A42A9A51547F8",
INIT_0B => X"1158936D20601A98A10200308A002E240010BFC0600002AFFBE249420555A2A2",
INIT_0C => X"1A3401A3401A3401A3401A3401A9A00D1A00C000850400A11414C005005000B5",
INIT_0D => X"10080C60AB0F42A8046282000DBFFF13D059280201948B029029409A3401A340",
INIT_0E => X"6FFFF8000F8F80281A16A1504302058102C0816244B82A0CA25907D0AA015874",
INIT_0F => X"0080A40000283D80000001402000283D80000001402010901A7D694494192200",
INIT_10 => X"0000034000283D80000001402000283D80000001402002010000A00000000000",
INIT_11 => X"C000000000000081600002080341C00000000000008C00000410085380000000",
INIT_12 => X"81000006809076B2000040400001080581000000000000004810020002010000",
INIT_13 => X"1051620000003410040004080000000040026C00008828B10000001A00210909",
INIT_14 => X"00503A000000000042AC00044000228A8000000000801204212130400000D001",
INIT_15 => X"1000000001064180000000000010C02C000440000240000000000105B0001040",
INIT_16 => X"964C4A44A0C689FF3F9FFEC5D6DBFE0020096528A0B000000CC043EC60780008",
INIT_17 => X"6058160581605816058160581605816058160581605816058160581605816258",
INIT_18 => X"0581605816058160581605816058160581605816058160581605816058160581",
INIT_19 => X"17FFFFFFFFFFFFFFFFE058160581605816058160581605816058160581605816",
INIT_1A => X"AEBAEBFFF7FEFCFDF7FFFFFF5DE7CFCB773FFEFBFF3C7E1E779FFEFFF5060030",
INIT_1B => X"F7FBFDFEFF7FBFDFEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEB",
INIT_1C => X"000FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEF",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9E79E7BAF7DEBAFAFEFBEFBFFBFFDFFF7FCFF0FBFFDFF7EFDDFFFEFFE8000000",
INIT_1B => X"7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"0003F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"1084B030000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"6DA986092050306382C05A1C900000001FAE89016387B2A38B5000D03FA1C0C2",
INIT_05 => X"C0FFC338FF008048240426200081F147F1FB7F289B81FB8003A396D20940C3DB",
INIT_06 => X"098000C51000910100006C00426FFC7C202060445F1F2572060FE82671C607E1",
INIT_07 => X"0001020400440C41C000617FC0003021259CFDB01BF00020C001FF8040009800",
INIT_08 => X"2000200008020000000820440000100220489020000020000000000000000044",
INIT_09 => X"8004800E3CF3E0B1118C31747F000B33820209206FC9E80000000000220FD1FF",
INIT_0A => X"000687C0044040424B39FB6073C0010048A20000047C1F804FBEF01BEE8027E3",
INIT_0B => X"204A608142002A440492530C401049020221BF861FF0C06C493C800580000000",
INIT_0C => X"04003040030400304003040030600182001821011DCCC31222730048620C4382",
INIT_0D => X"000802004815010008840800405FF864008880661874500E00E0030400304003",
INIT_0E => X"1FFE81FF880EA000400098200C04080204010200810020C180904240400340B4",
INIT_0F => X"0000040403C0800002000E800003C0800002000E8000100780C2C30830806202",
INIT_10 => X"EE00000003C0800002000E800003C0800002000E8000017A0040000010003E02",
INIT_11 => X"000400003D80000020400DD01000000020003B80000000801AE0200000100000",
INIT_12 => X"000384000006118A080428846A80000000002000780C800180000201017A0040",
INIT_13 => X"808000001C800001F80020000001F8000000280807404000000E400001D01000",
INIT_14 => X"10000000003E020000280808AB01000000000F600000003A020000007080000E",
INIT_15 => X"652075000000000080786800010000280808BA0040000000F8800000A02003B8",
INIT_16 => X"223010010308025410082404A015F0FFE003182701B420800280C80201A81000",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_19 => X"17FFFFFFFFFFFFFFFFC080200802008020080200802008020080200802008020",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000080040",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"88280C4C7B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"00160090920C04800904848262220277E05152B280780D407428E723C01E1400",
INIT_05 => X"0F001CC000890026105810941C5C06800E008057641E00473C40680D32330C00",
INIT_06 => X"82541A028D584E40CB0583CCA0100000161F84322000DA8C40F003C80030780E",
INIT_07 => X"BF70E1C3BBBB1138AF7F888025340C0888430047040FEE182CA00044BC5827C5",
INIT_08 => X"CAFC1F1F07F0FE1C94F65B11555EAFFC1C306758B24197ABCDA467F2C9CF9B32",
INIT_09 => X"4FFB4730000011420A61080800B6E0C464258094101606D5A47A2A2098B02000",
INIT_0A => X"446000304A0488111084048E082D0ED020119D35F900002FB00105C01036D800",
INIT_0B => X"1FA599581D3A9583C105A892112C04C0A898403120071501A6C32222068A3050",
INIT_0C => X"789E07A9E0789E07A9E0789E070CF0184F038850A21008E514845AB510D0106D",
INIT_0D => X"9A95E954868AD0E52273F4AC2180000808061C01C48B0F81380CE0F89E07A9E0",
INIT_0E => X"4001120055704FC4A1624487E2489024481224091282C4300942A19439481842",
INIT_0F => X"5D65C3E3F01F52FFC1E0013C1F801F52FFC1E0013C1F8090423D38A18E3B15C9",
INIT_10 => X"118796BE001F567FC1E0013C1F801F567FC1E0013C1F9085DFBF7E15C06101C5",
INIT_11 => X"7E30F00C0270F3751F1FD00FECBF7E25C0700463E17B2C7F811FD7ADECC381C0",
INIT_12 => X"4190626D6491063597F9177B956EF378D33E4030061341F077C571F8F885DFBF",
INIT_13 => X"7F328E3082636B2807FFD80FE00007E03F7207D3E03F9167184131B5C40FE647",
INIT_14 => X"EFA0CAE06101C53E3647D3F144FCDD22B81C0098E57D9081FCE8C8520C4DAE20",
INIT_15 => X"1ADF08DBF81846A540049707E0FE3307D3F141FFB45478040570EED41F4FE047",
INIT_16 => X"C189601208A1502B4AA5584B4068000019A80098120BCA4C617635C938574FF3",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"A800000000000000000902409024090240902409024090240902409024090240",
INIT_1A => X"08208208831042720EE38E38AAF9C4C704DAB63A6D58B3C10BAE8E789AA09424",
INIT_1B => X"7C3E1F0F87C3E1F0F82082082082082082082082082082082082082082082082",
INIT_1C => X"0003E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F8",
INIT_1D => X"0000000000000000000000000000000030F007FFFFFFFFFFFFFFFFFFFFFFF900",
INIT_1E => X"155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AEBDEBA0000000000000",
INIT_1F => X"7FD5545FF8000155087FC0155F7D168B55007BFDF45085168ABA002E82145085",
INIT_20 => X"55568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D7FFFE1000554214555",
INIT_21 => X"FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF7FFC00100800175555",
INIT_22 => X"0002E974BA5D5168A00A2D142155005142010FFAE820AAFF842AABAA2AE95545",
INIT_23 => X"AAFF803FFFF5D2A821550000000BA007FD55FF5D7FC0145007FD740055041541",
INIT_24 => X"FFF082EBDF455D5142000082E82145FFD17DFEFFFD168BFFF780000BA007FE8A",
INIT_25 => X"FE3F000000000000000000000000000000000000000000000AAFBEAA00007BFD",
INIT_26 => X"6F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEBDFD75D2AA8A80EA8E2",
INIT_27 => X"1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B68B551475FAF6D1C55",
INIT_28 => X"7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA0000542A0070071C50BAFEF",
INIT_29 => X"B8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A8010E004924874825D",
INIT_2A => X"EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0120155EA568E870BAE",
INIT_2B => X"7ABA497A82FFAFD2A82485FD2415A105C21451ED42A002545E055FFBE81D0BE8",
INIT_2C => X"00B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6A5C7E3DFFFE90B45B4",
INIT_2D => X"F45592E88A0AFE80A8B0A0000000000000000000000000000000000000000000",
INIT_2E => X"A1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE975EFAAAAB5E1AF3AABF",
INIT_2F => X"1CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB65F520EBE9EF67D7BE",
INIT_30 => X"034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EBC11472800752117082",
INIT_31 => X"968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F3142341D5DEEBEF55080",
INIT_32 => X"7D58AC448B69C30E02116220415A9540AA854140A0A2047F353AAF6C77F7F20D",
INIT_33 => X"56EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7C91565455C141E4188",
INIT_34 => X"F0000001FF0000001FF01EABC4B8014174FF7DA80F52FEDE6BE93172D7D625B5",
INIT_35 => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F",
INIT_36 => X"0000000000000000000000000000000000001FF0000001FF0000001FF0000001",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000100000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"CA1800080848B0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000010822C00803804000001999EF9C00040B0002000001000640200001018",
INIT_05 => X"08000000000100030008010468220A0004000000001000032000200002100800",
INIT_06 => X"8201961000060444010081002080000080820100000008004880000000284000",
INIT_07 => X"210C18306788C0089409800001140082000100010405000410A0000010082500",
INIT_08 => X"0A48903121780004C6000311555521F183060AC564BF818B5EDFDE0044600301",
INIT_09 => X"45B103200000140802234800000584000004808400020011A4581A2200002000",
INIT_0A => X"021000000800810400000402083000510000050020820036200005C00026C000",
INIT_0B => X"40000002000A008182200000002404400000000000010500008020A022220040",
INIT_0C => X"68064680646A0646A06468064690321503234204020018200404010784700404",
INIT_0D => X"C417C16004C0B838221090240180000801000C8800000190191064620646A064",
INIT_0E => X"6000000010200200802100022008100408020401020040100142200E0E08A20B",
INIT_0F => X"0021E300B000000781E00140018000000781E00140018000002430E30E0615C9",
INIT_10 => X"0000024E0000000781E00140018000000781E0014001908400005E11C0610000",
INIT_11 => X"3C30F00C000000155800D00000003E21C0700000000F00118000000468C381C0",
INIT_12 => X"40900004A400081401A0000004041218503E4030060000004804318008840000",
INIT_13 => X"01208C30800025200003D807E000000000725201600090461840001340002606",
INIT_14 => X"0F00C0E06100000012D2005100409520381C00000005920004C0C81200009A00",
INIT_15 => X"00120850B8180625400400000010711200510004B41478040000005548016000",
INIT_16 => X"40002002080000000804000A0000000011A000100208C008611430A000040250",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"0800000000000000000100401004010040100401004010040100401004010040",
INIT_1A => X"8A28A2AC8090C69606492492C09945235D5F7E2A5040B80E1C863A2958000500",
INIT_1B => X"DD6EB75BADD6EB75BAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A2",
INIT_1C => X"0002E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BA",
INIT_1D => X"00000000000000000000000000000000C0FFFFFFFFFFFFFFFFFFFFFFFFFFFC00",
INIT_1E => X"FE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5555550000000000000",
INIT_1F => X"D1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7AEBDF455D2EAABEFF7F",
INIT_20 => X"5000015500557DF45AAD1400BAA2AE801550051555EFF7AA95400552AAAABAFF",
INIT_21 => X"F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB5500517DF555D2EAAA105",
INIT_22 => X"5552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBAFFD540155557FD5400",
INIT_23 => X"10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAABAFF842ABEF5D517DF5",
INIT_24 => X"E105D2E954BAF7AE80010082A97410557FEABFFAAFBE8BEFAAD1575EF557FFFE",
INIT_25 => X"056A0000000000000000000000000000000000000000000005D7FFDF4500043F",
INIT_26 => X"BDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC51C7A2FBD5490BFD1C",
INIT_27 => X"4924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA974BAF7FFEFB45FFAA",
INIT_28 => X"DB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2080BEF495FC71D5412",
INIT_29 => X"FD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4002D082082AB8B6DBE",
INIT_2A => X"487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF78E021FF1471FDEAAF",
INIT_2B => X"FF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545A2DA3FB7DAAD4AAAAF",
INIT_2C => X"00547AB8F550A8010E00492487482FFFE82A85EBAE2FFC55554ADBD7A2FFC7BE",
INIT_2D => X"545AAFBF7400FBF9424F70000000000000000000000000000000000000000000",
INIT_2E => X"74AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E5400021EF005162BEF047FD5",
INIT_2F => X"225FF5843404547184164AA5D2EBEEB0A2D555410D3555714F8338AAAA1D0AE9",
INIT_30 => X"409000512AEABFFDF79DCBF755962010BDCBBC21455D7FEABEF75550ACBB7582",
INIT_31 => X"0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3FFEAAEB083BC1000FF8",
INIT_32 => X"BD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF801F8BA0C57740BDAA",
INIT_33 => X"DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF5D16BABAA3EBC3157A",
INIT_34 => X"0000000000000000000596EBEF55080034E0A592A4AD00FB863550229BCABEB7",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000100000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0812",
INIT_01 => X"A145A00810790848048044A54E404340404000720885800802000906E4910200",
INIT_02 => X"5C010802020408040C455850AA055254090541A111200A104A0000000908B510",
INIT_03 => X"182002200C00004485264A001214912803150020218808002440854288890550",
INIT_04 => X"210302048014100160806B08702010102722C9E0412200651102418214049492",
INIT_05 => X"88510910540008812C06010018204342A58A08011290A1120A81230240018DCA",
INIT_06 => X"47450000022480090000210002A54C282122040CC9082D530085224410AA4204",
INIT_07 => X"2101020423408900940C402A900011012D41D518044C10025000AA8A50043D00",
INIT_08 => X"214912534123010085008010141521F020409260000100A00004428808102010",
INIT_09 => X"519D12041551589141A539C42A4C9608080004801700D10100311820A848E0AA",
INIT_0A => X"0244C28C000002025A81AE3048321002A700200900160AE42CAA839AA90442C1",
INIT_0B => X"42300225604004D080251121D0000400880178044355940A498C400004A00545",
INIT_0C => X"4F240472404F240472404D240441200692022B41365E53340EC6940564D012D6",
INIT_0D => X"00000620500403080A919000038AD03001C5080D1108C1009001404524045240",
INIT_0E => X"02AA40AA902408000010002220040C000201030201200C818098402082020438",
INIT_0F => X"0080A0000140000002000140200A8000000200014020100280E469C698353000",
INIT_10 => X"000003400A800000020001402009400000020001402008700000000010000000",
INIT_11 => X"0004000000000081400004C00000000020000000008C000010A0000000100000",
INIT_12 => X"0000000680004188000400840080000000002000000000004810000001420000",
INIT_13 => X"0000000000003409280000000000000040025000030000000000001A05100000",
INIT_14 => X"000000000000000042900000A100000000000000008012A2000000000000D026",
INIT_15 => X"4420300000000000000000000010C010000098000000000000000105400002A0",
INIT_16 => X"126000808200505448342228120090554000E00000000000088000A000000000",
INIT_17 => X"004010040300C0300C0300C0100401004010040300C0300C0300C01004010240",
INIT_18 => X"0400004000040000C0200C0200C0200400004000040300C0300C0300C0100401",
INIT_19 => X"9FC0FC0FC1F81F81F800C0200C0200C0200400004000040000C0200C0200C020",
INIT_1A => X"0410411823A4301040B2CB2CBACB002009C6B860185AA1491B0E2863E8001100",
INIT_1B => X"4A25128944A25128941041041041041041041041041041041041041041041041",
INIT_1C => X"03F25128944A25128944A25128944A25128944A25128944A25128944A2512894",
INIT_1D => X"00000000000000000000000000000000F0F007FFFFFFFFFFFFFFFFFFFFFFFC07",
INIT_1E => X"415410AA8415555087BFFF55A2AA800BAFFAE9540008002AA000000000000000",
INIT_1F => X"FBEAABA5D7FE8B555551421455D0002145552EBFEBA007FC21EFA2FFD75EFAA8",
INIT_20 => X"2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F784155EFA2AEBDEAAA2",
INIT_21 => X"5D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BAA",
INIT_22 => X"55D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AAAAAAAAAAAFFD157410",
INIT_23 => X"FFA2D17DFEFF7800215500557DF55AA80001FFAA80001550055575EFFF840215",
INIT_24 => X"0AA082EAAB5500517DF555D042AA10A284154005D0015410085568A00FF80175",
INIT_25 => X"8A2A0000000000000000000000000000000000000000000005D00020AAAA8002",
INIT_26 => X"C51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA800AAFFAA9543A08003",
INIT_27 => X"0105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF49040017D5D20B8EAA007F",
INIT_28 => X"A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492AA8BC7EBDFEAFEFFD0",
INIT_29 => X"6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6FFEFB6D555578F7DB6",
INIT_2A => X"0155C51D0092A071555D5E3AE821D00001FF0871C016DBED1FDE90E3A497492B",
INIT_2B => X"8007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6DBE8F401D7B6A000147",
INIT_2C => X"00410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C5BE8555400550A3842",
INIT_2D => X"0AAF7AA954AA00042AAA20000000000000000000000000000000000000000000",
INIT_2E => X"21EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE975EF005560B55F7AA80",
INIT_2F => X"A8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BEABEF057D68F5F5A000",
INIT_30 => X"BFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D57DF55D7AABFF5428AC",
INIT_31 => X"D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002CA8AA80800020AAF7F",
INIT_32 => X"680800FFF7AAA155F595542455512A975455D3AA8A005500151FF0C57401E5F3",
INIT_33 => X"7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A2AA801455D7FE8BFFF",
INIT_34 => X"00000000000000000000C3BC1000FF8409000512AEABFF5D79FCAF774AE005BE",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000200000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380206",
INIT_01 => X"014C9A40408001683C0462C99E004B61404040028804A0080A000D16A0990A0C",
INIT_02 => X"4809A902031800444460589C66E331352180D468B8240E600C0081110B80ACD0",
INIT_03 => X"DA14C2210C0001D235834A0648D60528330006810A80881068A80C029CC56330",
INIT_04 => X"20886819A02740ECD2107364B37569100A04C1E01CA52010990240420E205A08",
INIT_05 => X"5831803532410000260E272058232259954369000A506912018CA582480038D1",
INIT_06 => X"8381A014000200AC2190ED0002ACD99881822144C5A409430682800046294140",
INIT_07 => X"218408142740E2C0948C3066500071913209CC8004640102D003999552083D20",
INIT_08 => X"00409231296AA180C2000110001521F0810A92E7402F00AB0016CA080C600111",
INIT_09 => X"41B112014D30E43802A76DD09905882B010605A01A4941010211088A2A43A399",
INIT_0A => X"4A12D9820880832264119D004860900104002008000F399606BC07998BA546AC",
INIT_0B => X"42522013604080D084A01001C8302D00008153000731C3000988C0040A224110",
INIT_0C => X"602406824068240602406224068920151203030032545B7404D7804566594796",
INIT_0D => X"080600E04C442068088590000999C8E84041086C001091009001406824060240",
INIT_0E => X"E6660599902600209021204A010E1C850C428521C208480021D842081A03E231",
INIT_0F => X"0090000003200000000010002008A00000000010002008038666928B28A65300",
INIT_10 => X"000801000A200000000010002009E0000000001000200A380000000000000000",
INIT_11 => X"0000000000000088000002D00000000000000000028010001620000000000000",
INIT_12 => X"0000008201021C88000048800280000000000000000004000010000003600000",
INIT_13 => X"8000000000041019980000000000000040802000068000000000020805B00000",
INIT_14 => X"0000000000000000C020000C8300000000000000008200AE000000000010402B",
INIT_15 => X"41003100000000000000000002008020000C3800000000000000012080001298",
INIT_16 => X"737420C20A01405468360022201185CCE0128410820000008088021C40A00008",
INIT_17 => X"2108721085218852188521885218852188521887210872108721087210872308",
INIT_18 => X"1086214872108621C852188421C852188421C852188721087210872108721087",
INIT_19 => X"26AA555AAB554AAB5561C852188421C852188421C85218842148721086214872",
INIT_1A => X"0410412881D0B0000092492480A981E063C638321450A08899A62C314A810508",
INIT_1B => X"EA753A9D4EA753A9D49249249249249249249249249249249249249241041041",
INIT_1C => X"BC4351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A9D4",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF82A",
INIT_1E => X"02AA00AA843DF55FFAA955EFA2D168B55557BEAA000055420000000000000000",
INIT_1F => X"5568A00087BE8BFFA2D155410AA8415555087BFFF55A2AA800BAFFAE95545080",
INIT_20 => X"D0002145552ABFEBA007FC21EF007FD75FFAA841541008002AB55AAAA955EF00",
INIT_21 => X"5D7FC0155005168B455D042AB45F7FFD741000042AA10AAAABFF5508003FF555",
INIT_22 => X"A5D7FC2010A2D1575FFF7AA975555D2E80145F78415545082EBDEAAA2FBEAABA",
INIT_23 => X"FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABFFF7FBEAB55F7AABDEB",
INIT_24 => X"B5555557DF55A2AEBDF555D2E954BA002EAAABA002A821EF5555554AA087BC01",
INIT_25 => X"203A000000000000000000000000000000000000000000000082E820BAA2FBEA",
INIT_26 => X"800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6FB7D5D7FEAA3808554",
INIT_27 => X"E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E1557D1475FAF45BEAA",
INIT_28 => X"AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2FBD55D7BE80004AA1E8",
INIT_29 => X"C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FFF5D0438140E2FA38B6",
INIT_2A => X"EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75D0A901FFFF801557D1",
INIT_2B => X"74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB455D20BDE00EBAAA8BC7",
INIT_2C => X"001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125FF002EADA921420871D",
INIT_2D => X"FFF5D7FEAABA0051400A20000000000000000000000000000000000000000000",
INIT_2E => X"75EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAAB55A28408145AAFFFF",
INIT_2F => X"D7145FBB8020A35D2ABEF55F7800015F087FEAA00007FEAB55FAD568AA2AFAE9",
INIT_30 => X"5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF55042AAAA007FD55558A7B",
INIT_31 => X"040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057968F575D003FF55F7D",
INIT_32 => X"52A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AAFFD5145FBAC9755F05",
INIT_33 => X"052ABFE10550415557085540000005156155FE90A8F5C082E974AAF7D57DF455",
INIT_34 => X"00000000000000000005500020AAF7FBFFFEF04552ABFFFF843FFE77C80825BC",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000100000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804002061080A284201081034809800A00230340007833522C82D04A16002",
INIT_01 => X"80439982183828490400050E12000340403008418984014902030106A0D10204",
INIT_02 => X"480108A000000000446418E01E80F00A41043118680402000800000009882390",
INIT_03 => X"0CA080210C0000408006480002001120260012603000000030808900888100F0",
INIT_04 => X"4403A609A055306B82C0705800CEE510082AC0A16B0350E3808041D03865D002",
INIT_05 => X"C0F20B36F0000901240626200820E26780E244A19A41E4020BAB06404001D312",
INIT_06 => X"434420151220118900806922406C3C7800201448DD9D2870020F228075A60715",
INIT_07 => X"2181000023480040840C001E180030032009700024641002C00187A440047C00",
INIT_08 => X"084830110160208004000001101121F220000260000100AA0004408000000001",
INIT_09 => X"519102063DF3E02B100B097407448F200A0209A041CA290102130C8800466478",
INIT_0A => X"8543D048006040064010E4007F62110105002002044007846124E0A00E0DC1EB",
INIT_0B => X"60020291404024808030512C40106D022203B1445810856A019400058F8404B5",
INIT_0C => X"052430D24305243052430D24304121A6921863013FD8807626EE000D64540284",
INIT_0D => X"28081080508104400A00800009B878680000880C1160410C90C143152430D243",
INIT_0E => X"81E0E18790012A00080102280800000202010102810020018098404110020004",
INIT_0F => X"0090000005E0200000001000200C6020000000100020000390E6C30830806204",
INIT_10 => X"000801000D20200000001000200EE0200000001000200A6A2000800000000000",
INIT_11 => X"8000000000000088000003B00100000000000000028000002EA0001000000000",
INIT_12 => X"80000082000251D80000C0044280000100000000000004000010000003282000",
INIT_13 => X"00002000000410121800040000000000408030000B8000100000020806F00000",
INIT_14 => X"0000100000000000C030000C9000008000000000008200FC000010000010403B",
INIT_15 => X"A500100000000100000000000200803000042E000200000000000120C0001590",
INIT_16 => X"30000800002400044934040AA231B63C20530801000410009889821040A00008",
INIT_17 => X"00401008000040300800004010000200C01000020040100802004030000002C0",
INIT_18 => X"000000C0300401008000000200C0100C01000020080000C030000000C0100802",
INIT_19 => X"325930C9A6CB261934C000200800004030040300800000020040100C03000000",
INIT_1A => X"8A28A2BD30264686668A28A2605145031C03F028000A1C2ED7831A2820244140",
INIT_1B => X"8D46A351A8D46A351AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A2",
INIT_1C => X"CFB068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D068351A",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF82B",
INIT_1E => X"54200000557FE10FFFBEAA10007FD7410FFAA97555082A800AA0000000000000",
INIT_1F => X"043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D168B55557BEAB45005",
INIT_20 => X"A8415555087BFFF55A2AA800BAFFAE9555508002AA000055574105D2A800AA00",
INIT_21 => X"087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAAA",
INIT_22 => X"0F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55A2AA955EF005568A00",
INIT_23 => X"AAA2FBD54BA080002145552ABFEAA007FC21EF007FD75FFAA8417410A2D14000",
INIT_24 => X"41000042AA10AAAABFF5508003FF55F7D568A00552EA8BEFA2AABDEAA087BEAA",
INIT_25 => X"50B800000000000000000000000000000000000000000000055042AB45F7FFD7",
INIT_26 => X"6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D5400F7A49057D08248",
INIT_27 => X"157428492E8008200043FE925571EFA380871C7028A28E3AF55F7A0925D7AADB",
INIT_28 => X"75C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA145",
INIT_29 => X"6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AAAEA8A9200249056D41",
INIT_2A => X"BE80004AAFEDB42028EBFBC2028BED152438AAA092492AAA4954281C0E2FB55B",
INIT_2B => X"FAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA007FC51C7007BD55D7",
INIT_2C => X"0041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEBAF7DF6AA00412EAABF",
INIT_2D => X"410FF84021EF0800154B20000000000000000000000000000000000000000000",
INIT_2E => X"AB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568A00FFFFEAA105D5155",
INIT_2F => X"955EF00042AAA25555410BA082E8201000043FE005D517DEBA0851574B2AAAEA",
INIT_30 => X"AAAA000804001FF005575408AA557FEB2FFAE975EF555168B55F7AA800BAF7AA",
INIT_31 => X"AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD568AA200557DE00AAA",
INIT_32 => X"07FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7D1550AAAA8002010F2",
INIT_33 => X"F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30800021EF55042AAAA0",
INIT_34 => X"000000000000000000008003FF55F7D5420BA5D2ABFEAAF7AEBDFF779A82AA43",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000200000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF0A0791B3FC1694378283C81FD996A091A32142007A336A20E03C040C002",
INIT_01 => X"A91FBDC4983088485C4A60000C24C26041280A00084000C8C212812EE2953231",
INIT_02 => X"C809AD5EB118E640A4F548FC011FF0002080000082ECC66609DB7DDDCB1FA036",
INIT_03 => X"4A120E4D3E4C90D294A31E824A52847A0B20640A88800000B8E0FD522885500E",
INIT_04 => X"001440849A2604001934800041110A71E2B068B110DB321C662AE22DC08A3448",
INIT_05 => X"370C14CA0E0800022446011C4E7F17907BEBD1AA65AE10571450DFC152522449",
INIT_06 => X"07319A109D129D450A846FE4E24C0305A1A5901C82416D05417118630839B88A",
INIT_07 => X"A5B56AD5A718C038AFFEA9FE39348C9204C389672407EE120EA5806E6C503AC5",
INIT_08 => X"C05896372728FF8C420619000003AFF4AD52A2C5D26F0EABCC96CD7AC4639902",
INIT_09 => X"5BD3571182080C000041080300F6F0C72221889C6FE20395A013282002B029F8",
INIT_0A => X"A23D203042444124098516CE0C2D13512410AD3CF8014005902DA6B2D1A4D810",
INIT_0B => X"645528937D5A85D3C4B0F883C10C24E0022B0E310612C2684CA16320A60A1185",
INIT_0C => X"288E3388E3208E3388E3288E330471904719C31438D04930ACE40FFD727C4304",
INIT_0D => X"8297A454544032252811E4AC2387F91008839C6CC413958D38C4E3208E3308E3",
INIT_0E => X"7FE0627FC25847C421516685844480204211200810028C38089AE00C894AA201",
INIT_0F => X"5D65E1E3C037E37FC3E0017C1F8037E37FC3E0017C1F900040261083080610CA",
INIT_10 => X"118796FE0037EA7FC3E0017C1F8037EA7FC3E0017C1F9300DFFFDE15D06101C5",
INIT_11 => X"BE34F00C0270F3754F1F8207FDBEBE25E0700463E17F3C7E054FF7BE6CD381C0",
INIT_12 => X"C090626DE40150459759573BBD6EF37D523E6030061341F07FC570F8FA00DFFF",
INIT_13 => X"6FE2AC3082636F301BFFFC07E00007E03F7263D383B7D1D6184131B7C1FEF64E",
INIT_14 => X"FFA0F0E06101C53E36E3D3EC84FDDDA8381C0098E57D923FDFC8D8120C4DBE0B",
INIT_15 => X"6FDF58DBF81C072540049707E0FE7323D3E43BFFF61478040570EED58F4F9397",
INIT_16 => X"00C108901822490448260224000040FC390250A2110B8ACC48B206A159A74FAB",
INIT_17 => X"08422080210882108C220842008821088230842208C20088210802308C2008C2",
INIT_18 => X"8422080230882108823080230842008C22084220842008C20080230802108C20",
INIT_19 => X"1092596D34924B2DA6884220842008821080230802108821084220842208C200",
INIT_1A => X"BEFBEFB7F7FE7EFEEE79E79EFAF2DDA73FBDCEDBFF9D3F0FDE0DB6DBF4208506",
INIT_1B => X"F77BBDDEEF77BBDDEEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"FED7BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF804",
INIT_1E => X"A800AAAAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF0000000000000",
INIT_1F => X"7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007FD7410FFAA97410082",
INIT_20 => X"A843DF55FFAA955EFA2D168B55557BEAB55005542000007FD74000055574BA5D",
INIT_21 => X"5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFFA",
INIT_22 => X"0F7D57FEBAFF80174BAAAD1555EF5555555550055574105D2A800AA00043FEBA",
INIT_23 => X"BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE95555080028A00A2FFFDE0",
INIT_24 => X"AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420BA5D2E821FFA2D5554",
INIT_25 => X"DFEF00000000000000000000000000000000000000000000000517FE10AAAAA8",
INIT_26 => X"D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC7010BEDF524AA5571F",
INIT_27 => X"1D74380851524BA5571D757DB6D5525EF555178F6D145178E00EBFBE8A101475",
INIT_28 => X"0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA147",
INIT_29 => X"92E8008200043FE925571EFA380871C7028B6AEBDF45B68A28B6DEBDF6DBEF1C",
INIT_2A => X"080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF55555057D1451524284",
INIT_2B => X"A552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45BEAA800AAFFAA9557D",
INIT_2C => X"0008517DE00AAAEA8A9200249056D4175C50920875FDA381C209256DFFDF420B",
INIT_2D => X"400F7FBC00BA55557DFF70000000000000000000000000000000000000000000",
INIT_2E => X"8A00AAFFEAA105D5155410FF84020AA0800154B2AAAA975FF5D7BC21EFF7FBD7",
INIT_2F => X"EABFF0051400A25551554BA0051400BA5551575EFF7D1401FF5D5568BE755556",
INIT_30 => X"AAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F78400145AAFFFFFEF5D7F",
INIT_31 => X"55421E75555400BA082E8201000043FE005D517DEBA0851574B2FFAABFF45FFA",
INIT_32 => X"7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF8002410FFD5575EF55",
INIT_33 => X"5D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7FFAE975EF555168B55F",
INIT_34 => X"000000000000000000000557DE00AAAAAAA000804001FF0055554088A557FEB2",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000C00000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000400322120040B313301C4389B2082",
INIT_01 => X"A74041CA38396849188160000C42424041000000090800090210090008110200",
INIT_02 => X"080108200C1000004465580000C0080100000000010432400800800009882050",
INIT_03 => X"080200010C234040842248600210812183806504488000103080014E88810000",
INIT_04 => X"0040504288A68210003120000000001002A0E8A910A072101000400A00203040",
INIT_05 => X"2800000400241801A52500094A02022014100128005004020010A1C044C02800",
INIT_06 => X"232000044084804914CA7C011AA3FC012122104CC0812D403280182308294000",
INIT_07 => X"2181020423488002940C0401D0480112000100004404004602447F8051223912",
INIT_08 => X"004812130160008304000000000021F020408264000108A00004400030400000",
INIT_09 => X"419102010104000A100348037F0584230A902A894008090343108802000FF407",
INIT_0A => X"B22D77C12052522400000400883011210000220006FC5FA400401484002447E0",
INIT_0B => X"60422291504420D084B0502044811428222300004611C57849A0150CA98A8561",
INIT_0C => X"1025B1025B0825B0825B1825B1112D8012D803003AD0413424E4014D627C0704",
INIT_0D => X"4404074040900B300A00810001A0021825E0886C0110916C96D15B0025B0025B",
INIT_0E => X"001E0800122100120499210A04A54652A12850962945180A14B44002CC020080",
INIT_0F => X"008ABA0030202100000001402068202100000001402067401026000000000031",
INIT_10 => X"00000341E8202800000001402068202800000001402062840000800000000000",
INIT_11 => X"8000000000000083D00052000100800000000000008CD0018400001200000000",
INIT_12 => X"800000069A48584000A0400000000005000000000000000048128D0002840000",
INIT_13 => X"80402000000034C1E000040000000000400FE000644000900000001A34000008",
INIT_14 => X"00003000000000004BA000112B0000880000000000807E80010010000000D1A4",
INIT_15 => X"0020250000040100000000000010CCE000198000020000000000010F80006028",
INIT_16 => X"0A728CA8C22540444924050CA9120603E0A2024048400010298432A002A00050",
INIT_17 => X"94E519465094A53946519425094A53946509425294E53946509425394E539625",
INIT_18 => X"425294E509425194E5294A519425094E5394A509465194A5294A519465094A52",
INIT_19 => X"3B1C618E38E38C31C71425294E53942519465294A53946509465394A50946519",
INIT_1A => X"8E38E39DB3B676F66EFBEFBEFAFBC5E73FC7F87A7D4ABFE7CFAFBE7BFA05004A",
INIT_1B => X"7F3F9FCFE7F3F9FCFE38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E3",
INIT_1C => X"6B23F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"00000000000000000000000000000000C0F007FFFFFFFFFFFFFFFFFFFFFFFC08",
INIT_1E => X"FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF0000000000000",
INIT_1F => X"AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFFBC0010AAD5574BA557",
INIT_20 => X"0557FE10FFFBEAA10007FD7410FFAA97400082A800AA08515555508043FE00F7",
INIT_21 => X"A2D5575EF55517FF55A2AA97400552AAAB45082E80155F7D1575EFFFAA955550",
INIT_22 => X"0FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD74000055574BA5D7FD7555",
INIT_23 => X"BAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000003DE1",
INIT_24 => X"B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE10AA803FE105D516AA",
INIT_25 => X"25FF000000000000000000000000000000000000000000000AAAEBDF45A28428",
INIT_26 => X"C7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49256DEB84104BAFFD15",
INIT_27 => X"B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE9756D145B401FFFFFF",
INIT_28 => X"DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A4904380824850381C5",
INIT_29 => X"851524BA5571D757DB6D5525EF555178F6DAAA495428412AAFB451C2A8017DE3",
INIT_2A => X"0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA2F1C50381471D74380",
INIT_2B => X"0A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D",
INIT_2C => X"00B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFFF1C7BD057D1C71FFE1",
INIT_2D => X"1FFAA84000AAFFD1401E70000000000000000000000000000000000000000000",
INIT_2E => X"75FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFDF55F78017400F78000",
INIT_2F => X"020AA0800154B2557FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2AAAA9",
INIT_30 => X"ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFFEAA105D5155410FF84",
INIT_31 => X"D5554B25551554BA0051400BA5551575EFF7D1401FF5D5568BE7AA80174AA082",
INIT_32 => X"AFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2AEA8A10082EA8BEFAA",
INIT_33 => X"557BC01EF55557DE00AA842AA0000516AABAFF8428BE7AAAEAAB55F78400145A",
INIT_34 => X"0000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000900000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0048201002842002C024500188000003000000003302300C018180006",
INIT_01 => X"020008402008404C042080000211024840000000080000080200010008110200",
INIT_02 => X"4801082248100000444008000080000041000000002222400800000009008010",
INIT_03 => X"0802010288A1484000020A400000002902006480088000003080040408810000",
INIT_04 => X"00004804890640004032030010000010008060E4100000140004500800403040",
INIT_05 => X"20000004004208016606010A0A20022000000000004000228010010080882000",
INIT_06 => X"030060004084004820906D311080020101000000008008011000000308290010",
INIT_07 => X"2100000023008002940C04000A4A010200018920646C10C50350002442003820",
INIT_08 => X"084812130160214204000000000121F000000244000100AA0004400920400000",
INIT_09 => X"419122810000081A00876882000590081100448A1000002350100CAA20002800",
INIT_0A => X"050280020100020400011640CC72602900044280028180242008069081244010",
INIT_0B => X"00200411508500B08805054C18024432A002400C99E410000080451100070014",
INIT_0C => X"05448054481544815448154481C22406A2406851201000200484950500F0145E",
INIT_0D => X"0144414A40000022880081511180036040044A013268E1205202480544805448",
INIT_0E => X"6000600010000020001102080102048102408120402800086098480008A20000",
INIT_0F => X"A2081210380021000001E003C0580021000001E003C042283426000000000021",
INIT_10 => X"00706801980028000001E003C0580028000001E003C044840000800009864038",
INIT_11 => X"80000330C00F0C0210807000010080000581C01C1C009201C000001200001607",
INIT_12 => X"8C2419101028D00020A2000000000005080082C180603A0E002A090404840000",
INIT_13 => X"8040204321188095F8000400061E001F800C202077C0009021908C4029F00008",
INIT_14 => X"00003009864038C10820201FAB000088026130071A00613E010011848322014F",
INIT_15 => X"6520350000640912058100F81C0108A0201FBA0002008239020F100880807BB8",
INIT_16 => X"114400C0002140144C2480200000040024A28400800044222980300CC4A0805C",
INIT_17 => X"2048120483204802008020082200812048120481200802008020081204812048",
INIT_18 => X"0880204812048020080200812048120080200802048320481204802008220080",
INIT_19 => X"2C208200010410400020C81200802008120C81204802008020C8120481200802",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000002A1050A",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"9840000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF818",
INIT_1E => X"5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04155550000000000000",
INIT_1F => X"AAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAAA97555F784174BAF7D",
INIT_20 => X"AAE955450055421FFFFFBC0010AAD5574BA557FFDFFF5555555EFAAFFFDFEFAA",
INIT_21 => X"A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00A",
INIT_22 => X"FA28000010552EBDE00007BEAAAAA2D14000008515555508043FE00F7AA97555",
INIT_23 => X"55557BD55FF00557FE10FFFBEAA10007FD7410FFAA97400082A800AAF7AE975F",
INIT_24 => X"B45082E80155F7D1575EFFFAA955555D51574AAAAFFD5545087FEAB455D516AB",
INIT_25 => X"7555000000000000000000000000000000000000000000000A2AA97400552AAA",
INIT_26 => X"9256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E1",
INIT_27 => X"B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7BFFF55FFA095482B6A4",
INIT_28 => X"2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF415",
INIT_29 => X"C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49003AFEFEBFBEAA001C",
INIT_2A => X"082485038F7A4905C7A28A070384120BDE100075EAA82BEDB470101C5B5057D1",
INIT_2B => X"5087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A101475D5400F7A490438",
INIT_2C => X"00AAA495428412AAFB451C2A8017DE3DF525FFFFA49756D495150492BEF1D255",
INIT_2D => X"A00555168A10002E9754D0000000000000000000000000000000000000000000",
INIT_2E => X"DF55F78017400F780001FFAA84000AAFFD1401E7FFAA97555A2AEA8A10AAD568",
INIT_2F => X"C00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215D557BF",
INIT_30 => X"028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7BC21EFF7FBD7400F7FB",
INIT_31 => X"FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2007FE8BFF080",
INIT_32 => X"D5155410FF84020AA0800154B2FF8402145A2AA954AA00043DE0000516AA10F7",
INIT_33 => X"005140000FFD140145007FE8BEF557BEAB55087FC215D555568A00AAFFEAA105",
INIT_34 => X"0000000000000000000AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"A140084000080048040100000202024040000000180800080200010048110204",
INIT_02 => X"080108020090000004655C000080000051000000002402400800000009008010",
INIT_03 => X"0002000100300C408422420002108108028065844880001030808D4288810000",
INIT_04 => X"0002584288A2C210003103001000001002A0E8C910A032541000090A00643040",
INIT_05 => X"2800080400645049A725010942220020140001A9005000004810A0C0044D2800",
INIT_06 => X"630400041404B141345A7C00426FFC01292214444081254102801A2308214004",
INIT_07 => X"21810204214080069408000008C3010200018920E06C0000021DFFA453263D32",
INIT_08 => X"084010110120018024000000000021F020408264000000080004400802400000",
INIT_09 => X"51B1004100040898128768820045142B0B902E895008080A1B13848A20002800",
INIT_0A => X"522920032052520400011641C460010D000000C8040100260008061081204010",
INIT_0B => X"4262229150012080102500211C81142880224000400411784920410C208514A4",
INIT_0C => X"0020000200002000020000200011000810008A55201000200484950004F0145E",
INIT_0D => X"40284301481509004885900101A0020964240109011890008011001020000200",
INIT_0E => X"0000200002210A320489000005A142D0A16850B6294D100A34B05242401340B4",
INIT_0F => X"00800008100001003C1FE00020080001003C1FE0002004401424008208041001",
INIT_10 => X"00000100080008003C1FE00020080008003C1FE000200080000001EA2F9EC000",
INIT_11 => X"01CB0FF3C000008000201000000081DA1F8FC0000080110080000002132C7E3F",
INIT_12 => X"3E6C00020040480040200000001004862CC19FCF81E000000010000200800000",
INIT_13 => X"004C11CF60001018000003F01FFE00004000000420800688E7B00008042000B8",
INIT_14 => X"000F251F9EC00000400004050002005D47E3F00000800084011607AD80004021",
INIT_15 => X"0000822406E5B85A3F830000000080000405000009AB87FB0000010000103000",
INIT_16 => X"1A768C68D260001448242704B912040002200640484000110104300042002018",
INIT_17 => X"B46D1B46D1B46D1B46D1B46D1B46D0B42D0B42D0B42D0B42D0B42D1B46D1B66D",
INIT_18 => X"46D1B42D0B42D0B42D0B42D1B46D1B46D1B46D1B42D0B42D0B42D0B42D0B42D0",
INIT_19 => X"200000000000000000346D1B46D1B46D0B42D0B42D0B42D0B46D1B46D1B46D1B",
INIT_1A => X"9E79E7B7F11E66C6FAD96D96520145052A1F5E2BD085122ED48F3AEB20840442",
INIT_1B => X"1F0F87C3E1F0F87C3E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"A6D4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF805",
INIT_1E => X"415555080000000087BEAA10F7803DE00FFAEBFFFF0800155FF0000000000000",
INIT_1F => X"80154105D7FC2145005155555F780155EFAAAEA8ABAAAFBFDE0055556AA005D0",
INIT_20 => X"87BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF552AA8AAA557FC0010F7",
INIT_21 => X"5D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF0",
INIT_22 => X"AAAAAA8B55F7D140010552E821EFAAAABDF555555555EFAAFFFDFEFAAAAAAB45",
INIT_23 => X"45557BE8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF5504000A",
INIT_24 => X"FFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F78402155AA8028A00A2D57FF",
INIT_25 => X"75D7000000000000000000000000000000000000000000000557BFDFFF55003D",
INIT_26 => X"FAE105D556AA10410E17555080E000280071E8A00EB8E3FE10F7AEBAFFF080A1",
INIT_27 => X"EA8AAA5571C2000FF8A17400557FC015514555757DFF8E175C7A2AAAAA82A2F1",
INIT_28 => X"FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF492",
INIT_29 => X"AF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A38492ABDE10EBDF7AF6DE3",
INIT_2A => X"5571FDFEF550E00082B6A0AFB55F7D1420104124821D7AAA0BDF6D415B575D7A",
INIT_2B => X"DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FFFFFFC7010BEDF524AA",
INIT_2C => X"00497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA001C2EA8A00F7800017",
INIT_2D => X"E00F7AEAABEF082E955450000000000000000000000000000000000000000000",
INIT_2E => X"7555A2AEA8A10AAD568A00555168A10002E9754D082E820BA08556AA00AAAABF",
INIT_2F => X"000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC21555D51575EFFFAA9",
INIT_30 => X"ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F78017400F780001FFAA84",
INIT_31 => X"843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215DA2FFE8ABA082",
INIT_32 => X"7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FFD540000000402145AA",
INIT_33 => X"5D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10AAAA975FF5D7BC21EFF",
INIT_34 => X"0000000000000000000007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000400000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000006",
INIT_01 => X"000009801830084C182060000C104268413C0A61590001D90213C10008110200",
INIT_02 => X"680108200010000054400C000080000041000000010002400800800009082011",
INIT_03 => X"0008000004002040000200100000000042800504488000103081880008C00000",
INIT_04 => X"00005042802A82100010030018000010000040C0100040140080040800003100",
INIT_05 => X"2000200400245001012100006002082000000000004000002010000040002000",
INIT_06 => X"2320400004040040144A7D000180020101000009808000000800001008210000",
INIT_07 => X"6100000021808000940800001800010200018B20206C01020200002441223C12",
INIT_08 => X"184010110120000004000000000061F000000244000081180004400000400000",
INIT_09 => X"4111002100040010008528820005100000900280000001000550860020002800",
INIT_0A => X"0080200520B23204000116404470900100402000000100242048025481024010",
INIT_0B => X"400000115040008002200000048034000002000000010712000000800F08A505",
INIT_0C => X"0000410004000041000400004100020000208201000000200404840284500016",
INIT_0D => X"00000120040000080000900201A0021924600088000000100100041000410004",
INIT_0E => X"60002000120002121C99024A00A14650A328519428651900142000000200A008",
INIT_0F => X"0000A20010200900000001400008200900000001400000001424008208041001",
INIT_10 => X"000002400820090000000140000820090000000140000A800000000000000000",
INIT_11 => X"0000000000000001500012000200800000000000000C10008400080200000000",
INIT_12 => X"0000000480004800002040000001000400000000000000004800010002800000",
INIT_13 => X"8041000000002401F80000000000000000025000274020800000001205D00808",
INIT_14 => X"004020000000000002900009AB00200800000000000012BA010100000000902E",
INIT_15 => X"652035000104000000000000001040100009BA000000000000000005400023B8",
INIT_16 => X"19028CA8D06540144C26832A1B0004000020024048400000090032A000000010",
INIT_17 => X"9425094250942509425094250942509425094250942509425094251946519465",
INIT_18 => X"4250942509425094250942519465194651946519465194651946519465194651",
INIT_19 => X"0800000000000000001465194651946519465194651946519425094250942509",
INIT_1A => X"34D34D1285B080201C92410480AB9A26667A46F345448020082E1C712A054008",
INIT_1B => X"1A0D068341A0D06834514514514514514514514514514514514514514D34D34D",
INIT_1C => X"2B60D069349A0D068341A4D268341A4D268341A0D069349A0D069349A0D06834",
INIT_1D => X"0000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF829",
INIT_1E => X"0155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA0000000000000",
INIT_1F => X"FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F7803DE00FFAEBFFFF080",
INIT_20 => X"780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555087BFDE00A2FBD7400F7",
INIT_21 => X"5D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA10F",
INIT_22 => X"A5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA557FC0010F78015410",
INIT_23 => X"45002EAAABA087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF780154A",
INIT_24 => X"E00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAABAF7D17FEBAA2AEBDF",
INIT_25 => X"8A92000000000000000000000000000000000000000000000AAFFE8A00552EBF",
INIT_26 => X"3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E",
INIT_27 => X"1FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E000280071E8A00EB8E",
INIT_28 => X"5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D556AA10410E17555087",
INIT_29 => X"571C2000FF8A17400557FC015514555757D5D71E8BEF147BFAE82A2DB555C71C",
INIT_2A => X"FFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A2AEADA38492EA8AAA5",
INIT_2B => X"2FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482B6A49256DEB84104BA",
INIT_2C => X"00A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D7000400155FFFBEDA8",
INIT_2D => X"B55FFAABDFEFF7D16AA000000000000000000000000000000000000000000000",
INIT_2E => X"20BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568BEF080402000F7AAA8",
INIT_2F => X"68A10002E9754D00517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00082E8",
INIT_30 => X"FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AEA8A10AAD568A005551",
INIT_31 => X"AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D51575EF555568BEF5D7",
INIT_32 => X"780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AAAE800AA552A97400A2",
INIT_33 => X"080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE00557BFDF55F78017400F",
INIT_34 => X"0000000000000000000A2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000800000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A14009821830284D182060000C10426840000000080000080200080000510204",
INIT_02 => X"0801080200100000046558040080000041000000002402400800000009008010",
INIT_03 => X"00020201040000D0842242024210810802006400088000003080054288C10000",
INIT_04 => X"0000400088020000003020002000001002A0E881108032100002000800203040",
INIT_05 => X"200000040000004924040108022000201000012800400010001081C040402000",
INIT_06 => X"030040040404804100006D2002A002012120004CC08125410200082308290000",
INIT_07 => X"2181020421408000940820001800010200018920206C01020200002440003C00",
INIT_08 => X"084010110120018004000000000021F020408264000000080004400800400000",
INIT_09 => X"511110010100008210010802004404230A000888400809000010042002002800",
INIT_0A => X"0000200000C04204000116404460910100082000040100240000000000004010",
INIT_0B => X"0AE22291404020902005002010000420A0200000400414684920410420200000",
INIT_0C => X"1120001200012001120011200011000090008840221000240484110000F05044",
INIT_0D => X"000803004C150100088480000980020000050001011890008011000120011200",
INIT_0E => X"000060001000020010010248040200010000800241000008009042404003E0BC",
INIT_0F => X"0080A00010202800000001402008202800000001402000000026008208041001",
INIT_10 => X"0000034008202100000001402008202100000001402002800000800000000000",
INIT_11 => X"8000000000000081400012000300000000000000008C10008400081000000000",
INIT_12 => X"8000000680001040002040000001000100000000000000004810000002800000",
INIT_13 => X"0001200000003408000004000000000040027000200020100000001A00000800",
INIT_14 => X"004010000000000042B00001000020800000000000801200000110000000D000",
INIT_15 => X"0000000001000100000000000010C030000100000200000000000105C0002000",
INIT_16 => X"03700080022100404D26A42EA01004002022000080000000018032A000A00010",
INIT_17 => X"0040100401004010040100401004010040100401004010040100400000000200",
INIT_18 => X"0000000000000000000000010040100401004010040100401004010040100401",
INIT_19 => X"0800000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"8A28A28D532A0CCC2A28A28A7AA344854A07F069CB8930AFD6A1AAA902A14148",
INIT_1B => X"6532994CA6532994CA28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A2",
INIT_1C => X"CC772B94CA6532994CA6572B95CAE532994CA6532995CAE572B94CA6532994CA",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF831",
INIT_1E => X"FEAABA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE100000000000000",
INIT_1F => X"8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA803DFFFAA843DF45FFF",
INIT_20 => X"80000000087BEAA10F7803DE00FFAEBFFFF0800155FF00042AB55FFD168B55AA",
INIT_21 => X"A2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE100",
INIT_22 => X"05555555EFF7FBC0145F78028A00A2D142155087BFDE00A2FBD7400F7FBFDFFF",
INIT_23 => X"FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555007FD741",
INIT_24 => X"EAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB55AAD168ABA002A975",
INIT_25 => X"8E00000000000000000000000000000000000000000000000557BE8BEF007FFD",
INIT_26 => X"38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E071D7AAFBEFB455D71F",
INIT_27 => X"42AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1E8B6D002090482B68E",
INIT_28 => X"D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D7000",
INIT_29 => X"2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD5410490A3DFD7F7A4821D7A2",
INIT_2A => X"410E175550071D54104951555D7EBF5C5155E3842AA00BED1421450871FFE00A",
INIT_2B => X"5BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82A2F1FAE105D556AA10",
INIT_2C => X"005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A38410E2ABD749516FB5",
INIT_2D => X"555A2FBFDF455D556AA000000000000000000000000000000000000000000000",
INIT_2E => X"8BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC01EFA2FFD7545AAAE97",
INIT_2F => X"AABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D56",
INIT_30 => X"EBFF45F78400155A2D57FE00552EA8A00082E820BA08556AA00AAAABFE00F7AE",
INIT_31 => X"D54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00FFFBD5400082",
INIT_32 => X"AD568A00555168A10002E9754D085155410085557555AAD557555A2802AA10FF",
INIT_33 => X"002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAFFAA97555A2AEA8A10A",
INIT_34 => X"0000000000000000000555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000008FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400986B830284D1820E0000C3642484000000008000008820009080A512220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"00080D4912E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"000048048002400048150300100002504230C8D9109032100020160880223000",
INIT_05 => X"220004440040080142020015001004A01200012840440000B01088C0005C2400",
INIT_06 => X"431018040014804920906C74B320020121210045408165445220082008211002",
INIT_07 => X"A5B1220421408004A56E840008B90D0200018B60A0650D450FC800644A0438A0",
INIT_08 => X"485816170760268E04000000000323F42C50826490640D28088445B0E0419003",
INIT_09 => X"41F1654100000818128728820024002B3B01AC9540080824CA13008820A02800",
INIT_0A => X"0000203600E06204000116C14474A3650048CE64E40100260048025481024810",
INIT_0B => X"08C32E915D9C208070042420180D24C8802000284007126A4D21262C20200404",
INIT_0C => X"31CA821CA831CA831CA821CA83165410E541085102000024040490A000D01056",
INIT_0D => X"812203360410110A4000840E3180021040465501011934A005101431CA821CA8",
INIT_0E => X"60006000101004A01811064B050204810240812241280D00200A08044290A088",
INIT_0F => X"482A01AAEC3602330CD2A02952DC3502330CB4A0318B41400024008208041011",
INIT_10 => X"0144C0155C3502330CD2A02952DC3602330CB4A0318B5600C587149B6D0141B0",
INIT_11 => X"083B6A51005956308D1E8202C436375908AA840AD4513437640F15245B455163",
INIT_12 => X"62F47B2872400044959BC42B1060F0D036B80B548523136C158878D8FE04E587",
INIT_13 => X"0A2699AAA3794392000D81852B0A050C224180062085134CD1719564E020C670",
INIT_14 => X"C50500D94C8121713C02B555101C90705D71009604140C0418CE0C378F0B2701",
INIT_15 => X"828E024D8C50965A40821568A06113801505010334AA73AA0666DAC20AD57400",
INIT_16 => X"123408C0822040544D248604B2100400100084008001D0113920060CDC06A27C",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"0080200802008020080200812048120481204812048120481204812048120481",
INIT_19 => X"0000000000000000002008020080200802008020080200802008020080200802",
INIT_1A => X"2082082815220A4A380000002A8313044020C0605885026853A1082100A00142",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000008208208",
INIT_1C => X"F070000000000000100800000000000000000004020000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF801",
INIT_1E => X"FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA0000000000000",
INIT_1F => X"2A801FFF7FFE8A10A28000000007FC2155F7D155545AA80001EFAAFBEAB45557",
INIT_20 => X"AFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2AEBFF45FFAEBFEAA00",
INIT_21 => X"FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEFA",
INIT_22 => X"5557FC2010002A80010A2842AAAA007BFFF4500042AB55FFD168B55AA8000010",
INIT_23 => X"EFFFD540000080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00557FF4",
INIT_24 => X"FEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021FF5D00154BAF7FBE8B",
INIT_25 => X"70AA000000000000000000000000000000000000000000000A2FFD741055003D",
INIT_26 => X"071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142ABDFC7F78E3FE28B6840",
INIT_27 => X"EBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007BC217DEBDB55555AA8E",
INIT_28 => X"AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92BEA",
INIT_29 => X"BDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA28A28BFF082ABAE10B6",
INIT_2A => X"080A175D708517DF7D497BC5028142A87000A28A2AA92007FF8F7D00042AB7DE",
INIT_2B => X"F5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00EB8E3FE10F7AEBAFFF",
INIT_2C => X"00B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E00B6DB6AA28A280001F",
INIT_2D => X"F55F7AABDEAAF784154BA0000000000000000000000000000000000000000000",
INIT_2E => X"01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBFFEF007BE8BFF5D2ABD",
INIT_2F => X"BDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BA087FC",
INIT_30 => X"AA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF080402000F7AAA8B55FFAA",
INIT_31 => X"7FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D5555FFAAA",
INIT_32 => X"AAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D2E95400A2AEA8A0000",
INIT_33 => X"FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA082E820BA08556AA00A",
INIT_34 => X"0000000000000000000FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000800000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702484000000008000008820009280A553231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"421A0A0012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"02004000890200001837830011998C31C09060DC104000102002140900003548",
INIT_05 => X"240000C400000001E404001F064000A00800000020480010A4100100001C2000",
INIT_06 => X"0300D800C1960C4400006E10B900020181840001008040057840001308212000",
INIT_07 => X"652428112180C03E8E5A2C800A3F018200418927E06686450FF8006460003A00",
INIT_08 => X"9840903525281D4F460409000000E3F08D1202C5C26A0719CC96CC7BF4629900",
INIT_09 => X"491175E10000041000C52882008600843001E09F0000002CF810200022302800",
INIT_0A => X"00002000030003040081164FC469227D2008CFE09A8180248009021091004810",
INIT_0B => X"00010C13499F01B33A00ACC0000F04F800000011800000000000433800000000",
INIT_0C => X"20CBC20CBC30CBC20CBC20CBC3065E1865E1000100000820040482B280504016",
INIT_0D => X"E7F3F01F40401C17E800C7FF3B80020000035780460124F16F06BC20CBC30CBC",
INIT_0E => X"00002200004005002001408400000000000000000000053A4096F80705FA0201",
INIT_0F => X"7B2C53F2FC16691DB587201EDDF4162B1DB527201EDDC46070241001000200F5",
INIT_10 => X"01D5CC9794162B1DB587201EDDF416691DB527201EDDD884272592D6246FC1B1",
INIT_11 => X"8E995D5A825DBA569F9FF02547068618CD3CC45B7863AE7EC00D4B122A67DF2A",
INIT_12 => X"CA5C33717461C045B5B182019473D19D7CCD856106F31A683621BDFC28800725",
INIT_13 => X"0A652CC8E3538BBA01624E51AA6C0469AC5493F5688532966471A9C5F6208C6C",
INIT_14 => X"41E1F5759001B4AA1853E6D5144AA9C914C8608D2724A4C4118D992B866E2FB1",
INIT_15 => X"825682D4A36C0B0B4B85112B2C4A05D3E6D5051893335EB0072AA85A4F9B7400",
INIT_16 => X"00800000082100544D248020000004001DC0800000010E7F70171401DE07EAD9",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0401004010040100401004000000000000000000000000000000000000000000",
INIT_19 => X"0800000000000000000040100401004010040100401004010040100401004010",
INIT_1A => X"249249120780800016A28A288028DCA30444409B054A88C5890486582A210108",
INIT_1B => X"32190C86432190C8641041041041041041041041041041041041041049249249",
INIT_1C => X"007592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2592C864",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF83E",
INIT_1E => X"0000AAAA843FE0008557DFFF0800020105D557FEAA00557DE100000000000000",
INIT_1F => X"AA8200000557DFFFF7AA80000082ABDF5508557DF45002ABDFFFF7803DE10AA8",
INIT_20 => X"07FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AAD5420000051555FFA2",
INIT_21 => X"F7FFE8A10A28000000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA0",
INIT_22 => X"05D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45FFAEBFEAA002A801FF",
INIT_23 => X"FFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA000028A1",
INIT_24 => X"BFF002ABDE00A2AABFE10082ABFFEF085542000000417555002A820AA08557DF",
INIT_25 => X"DE10000000000000000000000000000000000000000000000AAD155555A28428",
INIT_26 => X"BDFC7F78E3FE28B684070AABE803AE38145B78FD7000005010495B7AE921C517",
INIT_27 => X"547038145B505FFB6A487000005F7AFD7F7A482038002EBDF6D005B78F7D142A",
INIT_28 => X"2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00BED",
INIT_29 => X"BA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FFF1FDE821C003FE001C",
INIT_2A => X"F7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5D517DEAABEAEBFF7DE",
INIT_2B => X"5142082082005F7DFD7F7A482155BEF1E8B6D002090482B68E38FC7BE8A3DF7D",
INIT_2C => X"00B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FEF085F4703814001055",
INIT_2D => X"410007FEAA0055517DE000000000000000000000000000000000000000000000",
INIT_2E => X"FFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802AABA5D7FEAB45080015",
INIT_2F => X"FDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FEAB45F780020BA082EB",
INIT_30 => X"57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FFD7545AAAE97555A2FB",
INIT_31 => X"557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BAF7D1400BAFFD",
INIT_32 => X"7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA28428A105D7FEABEF55",
INIT_33 => X"087BD54AA550402145550000010087FFFF45F78402145F7D568BEF080402000F",
INIT_34 => X"0000000000000000000F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042604001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00020201926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"00104884880A4400403000004800027102A0E88110D83210642EA809C0203040",
INIT_05 => X"27000004004828032646000826080C201A008128044E00754010C9C192D82400",
INIT_06 => X"43000004080480492A946CE10320020121258044408125410270082308213800",
INIT_07 => X"A581424525408000AE2AA8002BC00D020003896020658FC4030000246E543AE5",
INIT_08 => X"4840101107200B80040210000002ABF02450A264002C80080004416800419000",
INIT_09 => X"4B531001000008001041080200B660E30B200C8840080A920651020002802800",
INIT_0A => X"0000203240E46204000516C04468C10100540034AC0100259001004010025010",
INIT_0B => X"04462E91440020905200A42209002420002800284002026A4D21758400000000",
INIT_0C => X"10000000000000010000000000000008000000000000002004040AA080504004",
INIT_0D => X"00000360401021280800E4000B800610C8410000A11210000000001000000000",
INIT_0E => X"6000600040D045E4195104D5854284A14250A12A512A8808289840084A020080",
INIT_0F => X"9E07A80948354B6E68982167061037496E683821670620681024000000000008",
INIT_10 => X"10B456587037496E689821670610354B6E6838216706220431961CA985D48094",
INIT_11 => X"186A91674011CE61403562274AA49CD594CF00039C7C414B6509DA22652138E5",
INIT_12 => X"3014780CC8604040424A5323845932E620295879818170304B2F5002C2043196",
INIT_13 => X"654B9104A328665603148895D44E0251142B42A3D8B2A5C8825194328A2E6A98",
INIT_14 => X"A6C6A465AA0091482382B17614F2202858EE300991415B45CD5306028F019451",
INIT_15 => X"08DC8047F17D1C7C3C02128E587D6A02B17605A130A4E8BF002258850AC5DC06",
INIT_16 => X"123508508220808048260604B2100C00022084809000D000393722A14000052E",
INIT_17 => X"284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A",
INIT_18 => X"84A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1",
INIT_19 => X"000000000000000000284A1284A1284A1284A1284A1284A1284A1284A1284A12",
INIT_1A => X"BAEBAEBFF6FEFEFEEEAAAAAAFBF7DDF77F9FBEFBFF9F3F0FDFCFBEFBF1228154",
INIT_1B => X"FD7EBF5FAFD7EBF5FAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAE",
INIT_1C => X"0077EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FA",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"57DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF0000000000000",
INIT_1F => X"7BEAB45552E80155AA802AB45AA843FE0008557DFFF0800020105D557FEAA005",
INIT_20 => X"82ABDF5508557DF45002ABDFFFF7803DE10AA80000AA087BD75EF087FFFFEF55",
INIT_21 => X"00557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAFFAE820AA5D55575550",
INIT_22 => X"FA2FBD7545FFD157555085140010F7AEAABFFAAD5420000051555FFA2AA82000",
INIT_23 => X"BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AAAEA8BF",
INIT_24 => X"EBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574BA557BE8A10A284154",
INIT_25 => X"ABD7000000000000000000000000000000000000000000000A2D155410F7FFFF",
INIT_26 => X"05010495B7AE921C517DE10A2DB50482147FFAF554971D0492E3F1C71C7BE8A2",
INIT_27 => X"1D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE803AE38145B78FD70000",
INIT_28 => X"A4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA1C7",
INIT_29 => X"45B505FFB6A487000005F7AFD7F7A482038AADF47092147FD257DFFD568A82FF",
INIT_2A => X"5D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000FFAAAFBFFBED5470381",
INIT_2B => X"24171EAA10B680124BAFFAAAFB45007BC217DEBDB55555AA8E071D7AAFBEFB45",
INIT_2C => X"00B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C20821C002AA92FFDF5748",
INIT_2D => X"010AAD157545F7AEA8B550000000000000000000000000000000000000000000",
INIT_2E => X"AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC00105D7BE8B55085142",
INIT_2F => X"BDEAAF784154BA5D5140145007BE8B55087BEAB555D04001EFF7AAA8B55F7802",
INIT_30 => X"FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007BE8BFF5D2ABDF55F7AA",
INIT_31 => X"AEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F780020BAA2FFD54105D7",
INIT_32 => X"AAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAAFBC0155085540000FF",
INIT_33 => X"5D042AA00F7FBD5410085568A10FF80020AAFFAABFF55087FC01EFA2FFD7545A",
INIT_34 => X"0000000000000000000F7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000CFFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"0002074F200904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000480488024000403000000000001002A0E881108032100002000800203040",
INIT_05 => X"200000040040080126060008020000201000012800400010001081C000402000",
INIT_06 => X"430000040004804920906C200220020121200044408125410200082308210000",
INIT_07 => X"A5A14285A15080008768A80008000D0200018B202067AF100A00002442043820",
INIT_08 => X"4850101105205380040000000000A7F42840A264920406080004400A00409002",
INIT_09 => X"411110010000080010010802000400230B000C88400808000211000002002800",
INIT_0A => X"0000203200E0620400011640446DA101004000002C0100240000000000004010",
INIT_0B => X"00422291400020900000002008002420002000004000026A4920410400000000",
INIT_0C => X"0000000000100000000000000100000000000000000000200404000000504004",
INIT_0D => X"0000022040100108080080000B80021040410000011010000000001000010000",
INIT_0E => X"0000600000000020181100400502048102408122412808082098400042020080",
INIT_0F => X"0040A100A42008000161C140000420080001C1C1400003201024000000000000",
INIT_10 => X"00022260042001000161C140000420010001C1C140001604E8084341CBA34048",
INIT_11 => X"2580E2B8802201014800C220A21829A302F1C024010C001124020C8C1A8A0396",
INIT_12 => X"0CA000048228404401004418012787124648157780120B8678C000801E04E808",
INIT_13 => X"072D04730000241000CB1325E78E0186030240000083B602398000120024ACA6",
INIT_14 => X"EF6F4163C480481506800004000CFD55196CB012481812049495C19400009001",
INIT_15 => X"800108B8FB61A0401200845594965000000400568D0CFB780055060500001001",
INIT_16 => X"123408408220000048240604B210040000008400800B0000090022A140068248",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"0481204812048120481204812048120481204812048120481204812048120481",
INIT_19 => X"0000000000000000002048120481204812048120481204812048120481204812",
INIT_1A => X"9E79E79FF3BEEEEEFE79E79EFAABCDA72E47F87BDF4EBAE7CFAFBEFB28200140",
INIT_1B => X"7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"FF83F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF83F",
INIT_1E => X"02ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA0000000000000",
INIT_1F => X"AE955455500155EF0804155EFAAD5554BA087FFFF55557BD54AAF7FBC01FFA28",
INIT_20 => X"A843FE0008557DFFF0800020105D557FEAA00557DE10A2AA801FFA28402000AA",
INIT_21 => X"552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400A",
INIT_22 => X"AA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF087FFFFEF557BEAB45",
INIT_23 => X"EF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA005568AB",
INIT_24 => X"555FFD168AAAFFAE820AA5D5557555002E80155A280000005D7FFDF4555517DF",
INIT_25 => X"0092000000000000000000000000000000000000000000000AAD1420AA087BD7",
INIT_26 => X"D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB4",
INIT_27 => X"E851FFB68402038AAAA955554900105FF0800175D7A2DB50482147FFAF554971",
INIT_28 => X"AAADB6D080A12410BE803AE38145B78FD7000005010495B7AE921C517DE10A2A",
INIT_29 => X"07FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2A0800BAE3F1C0092EB",
INIT_2A => X"B684070AA00516DABAA28402038B6803DE82F7F5D5410A2D568BC71C71D25D70",
INIT_2B => X"05D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D142ABDFC7F78E3FE28",
INIT_2C => X"00AADF47092147FD257DFFD568A82FFA4870BA555F5056D002A80155B6800001",
INIT_2D => X"145002AA8AAAAAFFC20000000000000000000000000000000000000000000000",
INIT_2E => X"00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFFF55FF84000AAAAFBC0",
INIT_2F => X"EAA0055517DE00A2AA955FFFF80020BAAAAA975450800001EF080417555A2FFC",
INIT_30 => X"0020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7FEAB45080015410007F",
INIT_31 => X"D56AB455D5140145007BE8B55087BEAB555D04001EFF7AAA8B555D557FE00A28",
INIT_32 => X"D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF803DE00FFD557400AA",
INIT_33 => X"082A80145F780020105D7BEAB45557BE8B45082EBFEBA082EBFFEF007BE8BFF5",
INIT_34 => X"0000000000000000000A2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000100000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"000440009282000001100000000000100220C8811080321000000228002A3000",
INIT_05 => X"200014C40000000100000000005C04A01000012A64400000145080C000422000",
INIT_06 => X"031042040804804100006EE4032002012120005540812540020008600831000A",
INIT_07 => X"21912244A14080008408880008000D0200018920206563000200002440003800",
INIT_08 => X"48501415032000800406180000002DF024408264000000080004400000430800",
INIT_09 => X"411100110000000010010802000400230A000880400808000450200000B02800",
INIT_0A => X"0000203000C042040001164044608101000000007C0100240000000000005810",
INIT_0B => X"0042229140002080000000200000040000200000400000684920000400000000",
INIT_0C => X"1000010000000000000000000100000800008000000000200404000010500004",
INIT_0D => X"00000260001001280000C4000300020000000000011010000000001000010000",
INIT_0E => X"400060000000000010010040040000000000000201000000000000004A000080",
INIT_0F => X"0000000000202100000000000000202100000000000004600024000000000008",
INIT_10 => X"0000000000202800000000000000202800000000000002000000800000000000",
INIT_11 => X"8000000000000000000002000100800000000000000000000400001200000000",
INIT_12 => X"80000000006000400080C0000000000D08120280000000000000000002000000",
INIT_13 => X"0040200000000010000004020010000000000000008000900000000000200008",
INIT_14 => X"0000308801400000000000040000008822110000000000040100100000000001",
INIT_15 => X"0000000004840717050000000000000000040000020000000000000000001000",
INIT_16 => X"023000000220000048240404A010040000008000000000000000020C40000008",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000200140",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"1420BAFF8000010082A954BA00003DFEF085155400F78428BEF0000000000000",
INIT_1F => X"843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD",
INIT_20 => X"AD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7AE95555A2FBE8BEFA2",
INIT_21 => X"5500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABAA",
INIT_22 => X"AA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FFA28402000AAAE95545",
INIT_23 => X"BA5D0015545AA843FE0008557DFFF0800020105D557FEAA00557DE10F7D1574A",
INIT_24 => X"0BAFFFFC20BAF7AEA8B45080417400FFFFC2145080015400AA802AA00AAAE800",
INIT_25 => X"DBFF00000000000000000000000000000000000000000000000516AA00A2AE80",
INIT_26 => X"50555412AA8ABAAADB40092E38E070280024904AA1C0438FD7005150438F78A2",
INIT_27 => X"A9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FFEDB55B6A080038E3DB",
INIT_28 => X"FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7E3A",
INIT_29 => X"68402038AAAA955554900105FF0800175D7E3FFEFBD70000124AA557FFDE10A2",
INIT_2A => X"1C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA38410038E38A2AE851FFB",
INIT_2B => X"0BE8E28A10AAA085082550A1057DBE803AE38145B78FD7000005010495B7AE92",
INIT_2C => X"001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A12410FFF1C017D14041040",
INIT_2D => X"B550855400AAF7AEBDFEF0000000000000000000000000000000000000000000",
INIT_2E => X"FF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA974AA0800020BA550028",
INIT_2F => X"57545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EFA2FBF",
INIT_30 => X"4020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7BE8B55085142010AAD1",
INIT_31 => X"002AAAAA2AA955FFFF80020BAAAAA975450800001EF080417555AAFFFDF45080",
INIT_32 => X"80015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7D17DF45007FE8AAA08",
INIT_33 => X"FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF7802AABA5D7FEAB450",
INIT_34 => X"00000000000000000005D557FE00A280020BAAAD140000A2AEBFFEF082A82010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000C00000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"0202115002BB10080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"2FE962000017102918900948514522CE09200C0D590569398ADBF8CC1E50E480",
INIT_05 => X"F05EA11E5600006B0800000038814B72A15B71D412E0AFD9C2990DA56FF0B55A",
INIT_06 => X"0640044150C025A0000000901A054F2C0A8030140BCC0460050690A95C8383D0",
INIT_07 => X"288500102F85203E8010D0AA9BC4800015001219D0550077373CAA8040006800",
INIT_08 => X"2064193920A2004B51400001414091EAA14881C0002701881B120203B7A80120",
INIT_09 => X"0409A02D965965200100104F2B00822512000000231520A024400800000ACCAA",
INIT_0A => X"0004B240028000342A00002FE00A3A1F06E649C005514AC40C082050010222D9",
INIT_0B => X"000A448C0082024AE50064B44000000000002A296AA000604838001980000000",
INIT_0C => X"044000440004400044000440004200022000200014808A02004200E540480212",
INIT_0D => X"0A80A5C8000102ED00440630004AD32400004000D58460018F6D3D8440004400",
INIT_0E => X"12AA28AA890BA00000024800480000000000000200802151025062C0BB400014",
INIT_0F => X"54E11C596A64003195933741477264003195555B418687E35836020814004049",
INIT_10 => X"99CF47DCB264003195933741597264003195555B4198843940076D296D0031F5",
INIT_11 => X"58486A556489347FE5F409CBC1362510695B6288743123C95251852041CD50A4",
INIT_12 => X"EAE2992046EB70026486035600CEC45CBCA809654B48163CCC895E1E043D4007",
INIT_13 => X"3A242DEA151848302BFD6D522B10C7EC71F6C1DB071D1216E078C4C1B1C74424",
INIT_14 => X"DAAABC982BE22267A2E2E4F44AA1DC5E37400C9EE1B7B638E8849D23C383298E",
INIT_15 => X"015998B28654565A003F0068E35352C1CAE48BFBF3A6C9B7B286B4DA8B93D037",
INIT_16 => X"009000040A8000452110A8442040D655602A102A0027E2C42320284086E6A2EE",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"1451451E96F2FC3C34F3CF3C2AC688AA263486D3260E34C0C3A7B451B0200000",
INIT_1B => X"7A7D1E9F47A7D1E9F4D14D14D14D14D14D14D14D14D14D14D14D14D145145145",
INIT_1C => X"0007D3E9F4FA7D3E8F47A3D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F4",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA0000000000000",
INIT_1F => X"80175EF0004000BA552A821FFFF8000010082A954BA00003DFEF085155400F78",
INIT_20 => X"2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D2E975EFF7D568BFFFF",
INIT_21 => X"AA8015400FF84001EF0000020AA5D00154005D043FF45555540000082EAABFFA",
INIT_22 => X"F5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555A2FBE8BEFA2843DE00",
INIT_23 => X"FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF557BEABE",
INIT_24 => X"4AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16ABFFFFAABFEAAFF84001",
INIT_25 => X"2092000000000000000000000000000000000000000000000FFFBE8BFF080017",
INIT_26 => X"38FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC",
INIT_27 => X"0925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E070280024904AA1C04",
INIT_28 => X"51420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB40092492",
INIT_29 => X"2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA410A1240055003FF6D55",
INIT_2A => X"BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC7557FC00BAE3AA9257DA",
INIT_2B => X"7F7AABAEAAF780051C70824851D7A2DB50482147FFAF554971D0492E3F1C71C7",
INIT_2C => X"00E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AABA08249756DF7D168BC",
INIT_2D => X"FFF552AAAAAA007BC00000000000000000000000000000000000000000000000",
INIT_2E => X"74AA0800020BA550028B550855400AAF7AEBDFEF08516AB55A2D16ABEFFFFBFD",
INIT_2F => X"A8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D04020AA002A955EFAAAA9",
INIT_30 => X"E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84000AAAAFBC0145002A",
INIT_31 => X"7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EF0800174BA002",
INIT_32 => X"85142010AAD157545F7AEA8B5500557DF45552A82000007BD74AAF7AEBDF455D",
INIT_33 => X"0804155FFF7D568B55FFAAAAABAFF8415545000015555A2FFC00105D7BE8B550",
INIT_34 => X"0000000000000000000AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000400000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"5295B6957FCBE0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"6DE90201BF90102103AF158E805428249851BFB2C106592088DBF8400A5055C2",
INIT_05 => X"403DA038338041EE341036BF36812841A19B68F40A807ED9C18114956FF081DB",
INIT_06 => X"00A0E2D7D3EAFF15800100FBFB333C1CBC303163670497AFF00291B3C0E20150",
INIT_07 => X"51C581123AEE54DE8008B719E61C10BBA5DAAFA9DDA1194D51E067BB00000000",
INIT_08 => X"0320A9392083056C2270E004400091181168C4D14002A110C902481FC0B42124",
INIT_09 => X"C51DFFC40C30E5F0182D0950190C0810BE00E9A76E4C6FFBE4700000B3038067",
INIT_0A => X"F7BC81C003C001674BB55B5FBB4BB4F26A19F70027CE86F047BEF19B6D94C1C1",
INIT_0B => X"0018CFC7429F326B9E822FFC00074D5A0AB033A3F330802966F74BFF8FCFB1F1",
INIT_0C => X"3EF3D3EF3D3EF3D3EF3D3EF3D3EF9E9F79E9E00185C44B91BC1740B7605040BE",
INIT_0D => X"CFEB69FF7A5F5AFFCCA787743FE67C21800367A28FC1AAF5CF6F3D3EF3D3EF3D",
INIT_0E => X"F99FD0678B87A0003000D8D02E00000000000000040025D3C21463D6BFF252D4",
INIT_0F => X"221ABD9CA854DFDD64A67D42C0F054DFDD64667D42C063E57A8F7B4594BB02C9",
INIT_10 => X"AA504801F054DFDD64A67D42C0F054DFDD64667D42C07237DFE5865F6D2BF232",
INIT_11 => X"8EAE7F5AB50D0806A9A2E0DFFF47DEDC496DA3181A0CC71440F9FBC3EFBB5AED",
INIT_12 => X"C3FC95949AEFF556EF9C75E7DCF1EB1B6E6FCDC87CB35FC94B36AECF3A33DFE5",
INIT_13 => X"AF5B6AAAE594A4C0DBFDAD94AA669809809FEFAF4157ADB55572CA527056E9C9",
INIT_14 => X"33F32ADD543430808BABAF50E1A5EB4BAEA45A250202FE0ADD39387F92B29382",
INIT_15 => X"523E865D4B1293AB6B90BF2F0E30EDEFAFD0B3FBD72E9E90D20A003FBEBF41AE",
INIT_16 => X"02F840000BCE0B6F67B3F845E017C833F6AAC02B002A2EFF22D4073DE83FB669",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9A69A6A4624C3434C0EBAEBA21B9001804F6E62029749701020B88A7CC0C0060",
INIT_1B => X"0D46A341A0D46A341A69AEBA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A6",
INIT_1C => X"00046A351A8D46A351A8D46A351A8D46A351A8D068341A0D068341A0D068341A",
INIT_1D => X"0000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA0000000000000",
INIT_1F => X"7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD17FFFF552EBFE00007",
INIT_20 => X"F8000010082A954BA00003DFEF085155400F78428BEFAAD168A000004020AA5D",
INIT_21 => X"0004000BA552A821FF5D00020BA552A82000552A821555D7FEAB55FF80175EFF",
INIT_22 => X"5AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EFF7D568BFFFF80175EF",
INIT_23 => X"55A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFFFFFDF4",
INIT_24 => X"4005D043FF45555540000082EAABFF00516AA10552E820BA007FEABEF0055555",
INIT_25 => X"AE920000000000000000000000000000000000000000000000000020AA5D0015",
INIT_26 => X"7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7",
INIT_27 => X"16AA381C0A07082497FEFB6D1451471EF007BD04920871F8FC7E3D56AB6DBEDB",
INIT_28 => X"7BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005150438F78A2DBFFBED",
INIT_29 => X"7D16ABFFE38E175EF1400000BA412E871FF550A00092492A850105D2A8015541",
INIT_2A => X"AADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5D7BFAEBA4920925EFF",
INIT_2B => X"2007FEDBD700515556DA2DF50492A2FFEDB55B6A080038E3DB50555412AA8ABA",
INIT_2C => X"000804050BA410A1240055003FF6D5551420101C2EAFBD7145B6AA2849248708",
INIT_2D => X"B550000175EFFFFBEAA000000000000000000000000000000000000000000000",
INIT_2E => X"AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFDFEFF7FBFFF55A2D16A",
INIT_2F => X"400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF5551555EF087FC200008516",
INIT_30 => X"A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800020BA550028B550855",
INIT_31 => X"7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002A955EF5D2E80010002",
INIT_32 => X"AFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FFD1575FF5504175EF5D",
INIT_33 => X"557FE8AAA000415410007BFFF450051555EFA2FBC0000A2FBFFF55FF84000AAA",
INIT_34 => X"00000000000000000000800174BA002E820105D003DFEF5D51420005D2ABFF45",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000CFFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"080BA868803F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"42016B0C401F58495C900A4859552A611D9A640F5903B2388004004C08A06008",
INIT_05 => X"7008000E0E508C01C28640000801133060E0032801E0202000991B708280B501",
INIT_06 => X"560000000022229A60B048048120FF040000000002C44D620F0228454C838100",
INIT_07 => X"58800A001D4033A004904087F9E3901218050018024110D6771C1F90C2856828",
INIT_08 => X"3020A82929A807B3731021400058C020000A9729400D10100420480202AC2140",
INIT_09 => X"0419002D86184A01018030430700802541420440022030041A814A0080064C1F",
INIT_0A => X"0000F0CA8428642430080438408A510185A200000045C18C0E0000A0820500B9",
INIT_0B => X"311324AA2373088479105D044A1022000001835C0C30C2E21480349D00100202",
INIT_0C => X"000C2000C2000C2000C2000C2000610006100100180A8062026000DC425C0301",
INIT_0D => X"10108003C00021002046088B5001FB3650D89844703657083080C2800C2000C2",
INIT_0E => X"007E281F840C00284A17210001060D8306C18360C1380A0260CB980840080810",
INIT_0F => X"9BBEF8E50B041029075982BF3873041029079982BF39748AA0AC800014804032",
INIT_10 => X"79BFD7F7F3041029075982BF3E73041029079982BF3F632C5F96D3C11555D5D7",
INIT_11 => X"A595405FC7F1CFEBC7586C4100A53162B47FD7E39FFEECE1598702345156AEA4",
INIT_12 => X"FE037ACFB88083A99E06271BB0CA207DFDD5920057E0B001B0EBCC79932C5F96",
INIT_13 => X"2A002DD51B6F7FC4A411D1E8D44517F14EAFE36E55150016EA8DB73E39464006",
INIT_14 => X"C30351452A13D55CFFA76E928E3891F148B30399F5FB7F28C800DFA06F5DF5CA",
INIT_15 => X"57DFEAEF1005475F1D1F608819CF0EE76E12C824ADD9089715F25FAF9DB84953",
INIT_16 => X"34041A41A0000010180C02801680460FC900052FA10DC0006DA4881C110155AC",
INIT_17 => X"60D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8",
INIT_18 => X"0D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D83",
INIT_19 => X"00000000000000000020D8360D8360D8360D8360D8360D8360D8360D8360D836",
INIT_1A => X"8A28A2891182C8A82E0820825945DF675C0770B9E11807E54587BEF8B0000000",
INIT_1B => X"2552A954AA5128944AAAA28A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A2",
INIT_1C => X"000128944A25128944A25128944A25128944A25128944A25128944A25128944A",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E954000000000000000",
INIT_1F => X"D568B55080028B55002E82000087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD",
INIT_20 => X"87FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA087FFFFFFFFFBFDF45AA",
INIT_21 => X"0051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE000",
INIT_22 => X"00804154BA55042ABEF5D7FD75FFAAD540145AAD168A000004020AA5D7BE8B45",
INIT_23 => X"10557FD7545FF8000010082A954BA00003DFEF085155400F78428BEFAA800000",
INIT_24 => X"000552A821555D7FEAB55FF80175EF5D00020105D2A97400082E95555085168A",
INIT_25 => X"24280000000000000000000000000000000000000000000005D00020BA552A82",
INIT_26 => X"E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A9",
INIT_27 => X"FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147FFFFFFFFFBFDFC7EBF5",
INIT_28 => X"003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092087",
INIT_29 => X"C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AADF6DB7DE3F5FAFC708",
INIT_2A => X"F78A2DBFFA28407038140410492550A2ABC7497BD25FFAADF4516DBED16AA381",
INIT_2B => X"8002E9557D1C516FA28417BD5545E38E070280024904AA1C0438FD7005150438",
INIT_2C => X"00550A00092492A850105D2A80155417BEFB6DEB8E175FF5D0E0500049209742",
INIT_2D => X"FEF552E974AA082A820AA0000000000000000000000000000000000000000000",
INIT_2E => X"DFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFFFFFFFFFFDFEFF7FBFF",
INIT_2F => X"AAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AA557FF",
INIT_30 => X"FFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D16ABEFFFFBFDFFF552A",
INIT_31 => X"FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087FC2000FFD56AB45A2F",
INIT_32 => X"50028B550855400AAF7AEBDFEFA280154BA550400000552AA8B45087FC01EFA2",
INIT_33 => X"5D2E974000804154BA082A975EF5D517DEAA007BD5545AAAA974AA0800020BA5",
INIT_34 => X"00000000000000000005D2E80010002A954005D2A82155087FFFFEFAAAA975EF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000400000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000010228001000000000000000000024001620280000000000354200004008",
INIT_04 => X"00016200001310090090004840004152C7208802590000388000004C08006000",
INIT_05 => X"7008000E0200000000000000000100302000000000E02000009900000000B100",
INIT_06 => X"00000000000000100000000000001B040000000002C42010010200004C838100",
INIT_07 => X"E0050A040041593104004500480090080A011202201400204204018000000000",
INIT_08 => X"30E409080188000021A0000100004082A140102B4020109801A4CE0037100100",
INIT_09 => X"00000005861840000000004301000B000000000001C1C0000000000000020C01",
INIT_0A => X"0000B0C0000000101400040C0408100000000000004540800000000000000099",
INIT_0B => X"000010000800011000000000000000000000BC0007C00008092C800080000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"08000EC0000000000000000010004B2000000000000000000000000000000000",
INIT_0E => X"0006280180040000000000000000000000000000000000000000000000000001",
INIT_0F => X"4451B81A70AB3006BA0011400760AB3006BA0011400680F02096834820000000",
INIT_10 => X"04082248A0AB3006BA0011400160AB3006BA0011400084C780687DBA82800808",
INIT_11 => X"796E80A00802301BC0A7531EDD98E73B02800804620D030F873EB49F30B80112",
INIT_12 => X"0000002044F091A860700FF9198AA115D5DA37F7A80C8A3604001C0664C78068",
INIT_13 => X"51AC9000000000314E01F9F30198600631448410A2A8D64800000081B0A936B0",
INIT_14 => X"0303842281C80A23004411AD661891F15148A4420804241526D6000000000985",
INIT_15 => X"35F3D282000C6C5456C84850F61050C411AD6284FDA861682805A04A1046B2E0",
INIT_16 => X"00000000000000000000000000004600C0013800003088004202304366A4A9D3",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"86186186851046260A9A69A6039045DD1F863808633005010063A20C90000000",
INIT_1B => X"930984C26130984C261861861869A61861861861869A61861861861861861861",
INIT_1C => X"0000984C26130984C26130984C26130984C26130984C26130984C26130984D26",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BA0000000000000",
INIT_1F => X"FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082",
INIT_20 => X"87FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7FFFFFFFFFFFFFFFFF7",
INIT_21 => X"080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA0",
INIT_22 => X"FF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFFFFFBFDF45AAD568B55",
INIT_23 => X"00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AAF7FFFFFF",
INIT_24 => X"B55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB55A2FFFDFEF5D2EBFE",
INIT_25 => X"04AA000000000000000000000000000000000000000000000AAFFFDF45A2D16A",
INIT_26 => X"FDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA00001",
INIT_27 => X"FFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7FFFFFFFFFFFFFFFF7FB",
INIT_28 => X"00001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92EBF",
INIT_29 => X"3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7F1F8FD7AAD16AB4500",
INIT_2A => X"087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D000000010087FFDFC7E",
INIT_2B => X"DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6DBEDB7FFEF552AB8E38",
INIT_2C => X"00B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E284971F8FC7AAD56DB6",
INIT_2D => X"FEF552E954AA0004000AA0000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFFFFFFFFFFFFFFFFFFFD",
INIT_2F => X"175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00557FF",
INIT_30 => X"56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FBFFF55A2D16AB550000",
INIT_31 => X"0402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AAF7FBFDFEFF7D",
INIT_32 => X"FFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7FFFFFFF552AA8BEF08",
INIT_33 => X"08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA0008516AB55A2D16ABEFF",
INIT_34 => X"0000000000000000000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000800000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"0001E6000053300B00D0005800000000000000407B0004BB830004DC3D01E000",
INIT_05 => X"F0FF433EFE022001C81080001101F977E0201C409BE1F10623BB000A100CF300",
INIT_06 => X"0F00100002E22EB440012C809B2FFF7C8E8840155FDC0000010E40087D8787A1",
INIT_07 => X"3B800000000000000008407FC800B0000000100600040000C205FF91C000F800",
INIT_08 => X"28C0B0300020852000002101554021F000000000000000090492260200002000",
INIT_09 => X"00000007BEFBC010002008FF7F00000000010018A81000041C401000004FFDFF",
INIT_0A => X"0002B7C0000008000000200000200A0C004408C2007D5FC800000240001227FB",
INIT_0B => X"000000000000000000000000800800A400000000000000008000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000800080000000",
INIT_0D => X"001000000100000020000800101FFB6000000000000000000000000000000000",
INIT_0E => X"07FE29FF800C00000001002040000000000000020480002E42429C0000080000",
INIT_0F => X"4D4E180010040000400000001E60040000400000001E6010003C000000000030",
INIT_10 => X"000094B1E0040000400000001E60040000400000001E60804000000400000000",
INIT_11 => X"02000000000033628000100100000004000000006170C0008001000004000000",
INIT_12 => X"000000295810000000A100020614148002000000000004307CC3CC0000804000",
INIT_13 => X"2000000000014AC000120200000000003F0D800020100000000000A4B0020000",
INIT_14 => X"0C0C00000000002E2D000001006204040000000005786C004000000000052580",
INIT_15 => X"0A0C0939BEE1810080200000E0CE0EC000010020000000000000AE8A00002002",
INIT_16 => X"8040400400C08080000000000049F6FFC0100000000000008008008000400010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000200",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C30C320624C1090D0F3CF3CD038001801C10000804482A60D09008269020010",
INIT_1B => X"86432190C86432190CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C3",
INIT_1C => X"000432190C86432190C86432190C86432190C86432190C86432190C86432190C",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"4174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804020100000000000000",
INIT_1F => X"FFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA000",
INIT_20 => X"87FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFFFFF",
INIT_21 => X"552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA0",
INIT_22 => X"FFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFFFFFFFFFFFF7FBFDFFF",
INIT_23 => X"EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA007FFFFF",
INIT_24 => X"FEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDFEFF7D56AB450000021",
INIT_25 => X"5000000000000000000000000000000000000000000000000F7FFFFFFFFFFFFD",
INIT_26 => X"FFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA08000",
INIT_27 => X"FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428087",
INIT_29 => X"FFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFFFFFFFEFF7FBFFFFF55",
INIT_2A => X"B6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AABEDF6FABAEBFFFFFFFF",
INIT_2B => X"7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7EBF5E8B550000071EF",
INIT_2C => X"00FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AAA497FFFFFFF7FBF8FC",
INIT_2D => X"FFF5D2A954AA0800174100000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410A2FFF",
INIT_30 => X"BFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFFFDFEFF7FBFFFEF552E",
INIT_31 => X"FFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00AAFFFFFFFFFF",
INIT_32 => X"2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAAD16AB450804174AAFF",
INIT_33 => X"087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA557FFDFEFF7FBFFF55A",
INIT_34 => X"0000000000000000000F7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"1094EC681244819000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"0001E6000053300F01D4587800446194F49020107F0012BBC00202DC3823EA82",
INIT_05 => X"F0F807BFFE000120080002341881F3FFF012412A9FE1E01013BF09404050F300",
INIT_06 => X"08808210996035A000006EC2E04FFFFC0A0000101FFE4036450E08247F878703",
INIT_07 => X"003400812A156C002822987FC830F40134CC74D002016612DE87FFE004008040",
INIT_08 => X"02348D2D00080C0C53400044114000000D022640B42406808790055043A82824",
INIT_09 => X"080AC707FEFBC110008420F7FF388B70A20389346FE8000580200800008FDFFF",
INIT_0A => X"4636FFC00080013029811240444A82422A828C03BC7D7FC15025B1AB6E85A7FF",
INIT_0B => X"2019480E63180855A492712CC01C49C20201BFE45FF0C004041DA2218A8A3151",
INIT_0C => X"648A3648A3648A3648A3648A366451B2451B210018C241102068006C620C0388",
INIT_0D => X"80050094104431200090080C621FFBE0008A94641165448C80C103648A3648A3",
INIT_0E => X"9FFEADFF8050250010030165290008800440022201082401A002000C48000201",
INIT_0F => X"48A004A6C0D2820302C005A83480D1820302A009B02B101390C0CB2830816202",
INIT_10 => X"8904831400D1820302C005A83480D2820302A009B02B021A85C0941150013180",
INIT_11 => X"8834600024D052C1051E0B92D400360520202682C19024B6164E300448510140",
INIT_12 => X"4093E22A2012418A9D1D44ADD9E0F174103820101C0B8160D5516259FA1A85C0",
INIT_13 => X"8AA288209E615100280DA0052000C5006402000206C55144104D510CC1B0D640",
INIT_14 => X"D50020C04023033C52009144231D902818100C90058010361AC808126C88660D",
INIT_15 => X"2386454988140600C0181500A13E830011008B0374007000B4E0CD00024500A0",
INIT_16 => X"0224004002000000703804008001F7FFF01B982B01258088C008CC41198A1220",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"0000000000000000002008020080200802008020080200802008020080200802",
INIT_1A => X"BEFBEFBFF7FEFEFFFE79E79FFFF7CFF77FBFFEFBFF9F7E0FDF9EFEFBF0000000",
INIT_1B => X"FF7FBFDFEFF7FBFDFEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000100000000000000",
INIT_1F => X"FFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080",
INIT_20 => X"7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAF",
INIT_22 => X"FFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFFFFFFFFFFFFFFFFFFEF",
INIT_23 => X"AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFF",
INIT_24 => X"FFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFFFFFFFBFDFEF5D2A954",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA00000",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAF7F",
INIT_29 => X"FFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFFFFFFFFFFFFFFDFEF55",
INIT_2A => X"082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA002A95400087FFFFFFF",
INIT_2B => X"FF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA",
INIT_2C => X"00E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50BA557FFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0000020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAFFFFF",
INIT_30 => X"FFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E",
INIT_31 => X"2E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410087FFFFFFFFF",
INIT_32 => X"7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7FBFFFFF552E954BA00",
INIT_33 => X"5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA557FFFFFFFFFFFDFEFF",
INIT_34 => X"0000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"8632CA211E4491D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"24B000808800040439245B221373581F97B0A8D1040F92000F42000047A00E58",
INIT_05 => X"0107C4410008816B105036B4180C000811E9BF2844021B1004045E4249500449",
INIT_06 => X"0111C2D50A46AE45281502E4A2200081ADA0E054402365774611E047020008E0",
INIT_07 => X"80BD5AA4BF5C91F840C1710010344DB9A808FDFF3DE0313014A2007540401804",
INIT_08 => X"EA212D6D481ADF0CE47CA21544009007A64EBD64049D028B93D9561A48F60276",
INIT_09 => X"0E48D500400015805060040080A2A0F4A82381B4000A0905A0283800AA500200",
INIT_0A => X"4E700838460402635019FBFE7FCA13520F8AAD050402204090090319A5002004",
INIT_0B => X"040F4A944B1AA313C0022AA0011C0DC0002800134000000849BCC3240A8A7151",
INIT_0C => X"70AA070AA070AA070AA070AA072550385503800500001840000C80B410014088",
INIT_0D => X"0A9CA0D458D131652A154CAC6B600085080B14004D1594832824A070AA070AA0",
INIT_0E => X"C00044000A1EC1C44140D101A54280A14050A028500A84F02842A24C594A0687",
INIT_0F => X"59E0C4E6C256690581800F1C3E82562B0581200F1C3F08145602280402080448",
INIT_10 => X"AB8581B602562B0581800F1C3E8256690581200F1C3F1238473F121000613383",
INIT_11 => X"0E1050083750B3E4275F829547008600C030374361FA2CEE046D48122C438100",
INIT_12 => X"C012A66F61154C019511628756231018500C00203E138061565160782238473F",
INIT_13 => X"AA612C0096C37B00D1724801A0009C606D1221D104553096004B61BCC1128C4C",
INIT_14 => X"41E0F0600035842E7601C2C4AC68A98810080AA825A890225189980254CDE608",
INIT_15 => X"637E00D0A1080301401C390320188321C2C0B13890105800D520AF94870B012A",
INIT_16 => X"22F110111B281A54753AA004002601001918008C10912A4440B24E8B58234A89",
INIT_17 => X"0882208822088220882208822088220882208822088220882208822088220882",
INIT_18 => X"8020080200802008020080200802008020080200802208822088220882208822",
INIT_19 => X"8000000001FFFFFFFFC802008020080200802008020080200802008020080200",
INIT_1A => X"9E79E7BFF3FEFEBEEEFBEFBEFBEFDFEF7F47F8FBEF5EB7E6CFEFBEFBE8289144",
INIT_1B => X"7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"0003F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000000000000000000",
INIT_1F => X"FFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFF",
INIT_24 => X"FFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFFFFFFFFFFFFF552A974",
INIT_25 => X"0010000000000000000000000000000000000000000000000007FFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0804154BAF7FFFFFFFF",
INIT_2B => X"FFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA",
INIT_2C => X"00007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000AAA2FFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804000100000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A",
INIT_31 => X"04174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAF7FFFFFFFFFF",
INIT_32 => X"FFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E974AA08",
INIT_33 => X"AAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA2FFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"5886C0201A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"0005EE040057700F40D08078500000D9218020407F0000BB8018A2FC380BEAC2",
INIT_05 => X"F0F817FFFE400800020224000405F7FFE0124002FFE1E0C517FF09111212F300",
INIT_06 => X"400000409120338860900482404FFFFC000000001FFC0832050E00047F97870B",
INIT_07 => X"00246801C41C3E81E872C8FFE900FC31348EFDF03BE15E22DA07FF92C2041020",
INIT_08 => X"6220280D2B025988311AB14155421006891A1089F6E200000022C140068EB902",
INIT_09 => X"0002021FFEFBC80000000077FF184B03010004002FE1F2900201000000FFDFFF",
INIT_0A => X"0006FFEA002020626995FBE077430001E7320006F87D7FA84024B0225A890FFF",
INIT_0B => X"241C482B20400CC52492710CC80060020A81BFE41FF0C2060481200180000000",
INIT_0C => X"040430404304043040430404304021820218210018C24110A860006C620C0312",
INIT_0D => X"001002001804800000952800001FFBF040C088669070510C90C1430404304043",
INIT_0E => X"1FFEAFFF805025E00853B92588000400020001000020A8018008002000014030",
INIT_0F => X"148484054395E27E428002A4200397E07E422002A420100382FCC30832A16382",
INIT_10 => X"788417000397E07E428002A4200395E27E422002A420110A51C01C0590401486",
INIT_11 => X"1A2490040590C08120558C1759BE1C05A0400383808800DA1929F728641100C0",
INIT_12 => X"00136006000215EA0A4833A32C8832050028603050014031B3950000C90A51C0",
INIT_13 => X"658280009A2030108B14AC05C00112405222088B8332C140004D101800CE7200",
INIT_14 => X"B6808060201281004228996085F10020180C030880D11019CE4000026C00C006",
INIT_15 => X"49DC7143F01C04240030720641E0A028996483A17204680410A04104A2659196",
INIT_16 => X"1000080080000000000002001201F7FFC0011C2F81A48080CA32800A0108152A",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"0000000000000000000040100401004010040100401004010040100401004010",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080002010FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA08",
INIT_33 => X"F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"0000745C200801000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"0001E6000053300F00D0007810042140C00000407F0000BB800000DC3801EA00",
INIT_05 => X"F0F8033FFE000000000000000001F17FE01240009BE1E00003BF00000000F300",
INIT_06 => X"000000009120110020100002404FFFFC000000001FFC0000010E00007F878701",
INIT_07 => X"00102050840950002802C87FC800FCAA035400001B918600C207FF8000000000",
INIT_08 => X"6234AD280B02500063AC2840001610020408178B600C24000136496087300042",
INIT_09 => X"00000007FEFBC00000000077FF000B00000000002FE0000000000000000FDFFF",
INIT_0A => X"0006FFE80000015406A800003388000025000002387D7F804024B0224A8107FF",
INIT_0B => X"20502000200000400490510CC00040020201BF441FF0C0000000000180000000",
INIT_0C => X"040030400304003040030400304001820018210018C0411020600048620C0300",
INIT_0D => X"800B00000000000000000000001FFBE0008080641060400C00C0030400304003",
INIT_0E => X"1FFEADFF80002080000000208800000000000000000020018000000000000004",
INIT_0F => X"009181008024A00043601100210024A00043C0110020901382CCCB28B0806202",
INIT_10 => X"040A03080024A00043601100210024A00043C01100209240C840C201D0210840",
INIT_11 => X"A604E0080820009908008341B000A8212070082002890010068320860C920180",
INIT_12 => X"00800082041205EC00044C1ACB66C37542082030281E0580001012811A40C840",
INIT_13 => X"27A004300004103160DB3005E000618040C022000593D002180002090166B406",
INIT_14 => X"FF20406040084210C062000C2A2DDD00180C04504086002CD680C0100010480B",
INIT_15 => X"04295C98F80400008040CC0582169022000C2876C404780028500160880012BB",
INIT_16 => X"0000000000000000000000000001F7FFC001B823018F00880008805241060208",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9EF9EFB263CC3090CABAEBAFF96857757B73E6089966B9EF9D5A220CC8000000",
INIT_1B => X"0F0783C1E0F0783C1EFBEFBEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF",
INIT_1C => X"0000783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2010000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020100000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA00",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00004000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"4909E6093253306F82D0007C80000000080E01007F8020BBC00040DC3801EA00",
INIT_05 => X"F0F8033FFF0240012C1400080291F17FF01241009BE1E00203BF80800000F392",
INIT_06 => X"0DC00CC0992033A062116E82404FFFFC0E0801101FFC0000010E08A07FC78701",
INIT_07 => X"00000000000000002802C87FC800F8000000000019810600C207FFF3C410D841",
INIT_08 => X"E8002000080281000008A0000014100200081000000000080480AE0000002000",
INIT_09 => X"80040007FEFBE031018C31F7FFBAEBC0020008086FE0000100280800000FDFFF",
INIT_0A => X"0006FFF800C04000000000003300800005000032387D7FE94FBEF2B2CB8DA7FF",
INIT_0B => X"20100000200000400490D10EC00040220201BF441FF0C0600000000180000000",
INIT_0C => X"04003040030400304003040030400182001821001DCCC31222730A49620C0300",
INIT_0D => X"000000000000000000012800001FFBE0008080641062400C00C0030400304003",
INIT_0E => X"1FFEADFF805025C0304001E58906088304418222C108A009A090400000000000",
INIT_0F => X"00100100000480000200100000000480000200100000100380F0C30830A06302",
INIT_10 => X"0008000000048000020010000000048000020010000000004040000010000000",
INIT_11 => X"0004000000000008080000011000000020000000020000000001200000100000",
INIT_12 => X"000000800002018C010000020800000800122000000004004000008000004040",
INIT_13 => X"2080000000040000001020020000000000800200001040000000020000021000",
INIT_14 => X"1000008001000000800200000021000020100000000200004200000000100000",
INIT_15 => X"0008400000000605000000000200000200000020400000000000002008000002",
INIT_16 => X"226410410346010000000400A011F7FFE0031823010400800000800001840000",
INIT_17 => X"2088220882208822088220882208822088220882208822088220882208822288",
INIT_18 => X"0882208822088220882208822088220882208822088220882208822088220882",
INIT_19 => X"17FFFFFFFFFFFFFFFFE088220882208822088220882208822088220882208822",
INIT_1A => X"0492410A048029890AD34D35FDD144A50CB5462D14997BE09E760AED04040000",
INIT_1B => X"6231188C46231188C49249249249249249249249241041041041041041049241",
INIT_1C => X"000B158AC562B158AC562B158AC562B158AC562B158AC562B158AC562B1588C4",
INIT_1D => X"0000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"94A7B2B1450000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"6FEBEF5FEC737AFBC6F85FDEB220109E1FEFFFE3FBA7FDFB9BD301DC3FF5F0D2",
INIT_05 => X"F0FFEB3EFFF7FDED3FBFF6A84383F177F5FB7FF59BE1FF980BBBB7FE6D21F3DB",
INIT_06 => X"FBE564C71268F3BBF5FBFC2A427FFF7C3E3A74667FDDB7FB870FF30FFDEF87F5",
INIT_07 => X"3BC18306396FBEC14489737FDC00B13BB79DFDB83BF4112AF205FFBDD3AFB93A",
INIT_08 => X"21E4391909B381B0B1F8E041051831FA3068D77E000030021324620C0B9C2060",
INIT_09 => X"D13D980FBEFBEBF30B8D79FF7F451F33CFD60FE8FFFDF54003B1D4223B4FFDFF",
INIT_0A => X"B5AFF7CFACFAFE776F39FF7077E29D83CFAB300B017F5FFE6FBEF73BEFB967FB",
INIT_0B => X"737AF3FD62601EDC25B3533DCEB07F262213FFC67FF1C7FBFB5EC9478D5DA3A3",
INIT_0C => X"5E3035E3035E3035E3035E3035E981AF181AE315BDDCC3B336F7C548667D47B7",
INIT_0D => X"100C0E60FB9FC3A80EF69A004DFFFF7FF5F9A06E19F4DA0E80E903DE3035E303",
INIT_0E => X"7FFFF9FF8FAFAA3ADEBFB9726BAF5FD7AFEBD7F7EFFD7ACDB7F947F0EA035CF6",
INIT_0F => X"0080A40403E8BD8002000FC02003E8BD8002000FC02010979AFFE36C36B86702",
INIT_10 => X"EE00034003E8BD8002000FC02003E8BD8002000FC020037B0040A00010003E02",
INIT_11 => X"C00400003D80008160400FD81341C00020003B80008C00801EF0285380100000",
INIT_12 => X"81038406809677FA080468C46A81080581002000780C8001C8100201037B0040",
INIT_13 => X"90D162001C803411FC0024080001F80040026C0807C868B1000E401A01F11909",
INIT_14 => X"10503A00003E020042AC080CEB01228A80000F600080123E232130407080D00F",
INIT_15 => X"7520750001064180807868000110C02C080CFA0042400000F8800105B02013F8",
INIT_16 => X"FF7EFEEFF3EEC3FF7FBFFBCB7FFFFEFFE00BFF7FEBF420800EC0CBEE61F81008",
INIT_17 => X"F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F7FD",
INIT_18 => X"5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7",
INIT_19 => X"37FFFFFFFFFFFFFFFFF5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F",
INIT_1A => X"A61861BAF15EAA6AFC38E38EA3AD8ADE7A48F0B366429F434AA9FC376DAE4432",
INIT_1B => X"130984C26130984C261861861861861861861861861861861861861861869A69",
INIT_1C => X"0000984C26130984C26130984C26130984C26130984C26130984C26130984C26",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"1085B0B041000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"6FAB975B6470BAF386C87A9CB00000001FEF9F23E3A7BDE79B5101D23FB5C0C2",
INIT_05 => X"C8FFCB38FF35B44C25ADE72041A3F147F5FB7F759B91FB880BA3B6FE2921CBDB",
INIT_06 => X"B98420C71408D113956AFD0842FFFC7C3032646EFF1DB7FA868FE30EF1CE47E5",
INIT_07 => X"0041830600640C415004637FC4003021259CFDB01BF80028E001FF8251AB9D1A",
INIT_08 => X"200822020842203000082050000110023068D030000028200000008400000051",
INIT_09 => X"90A4880E3DF7E2FB0B8E717C7F411F3BC6D60B60FFDDE440018AC4AA3B0FD1FF",
INIT_0A => X"042787C5AC5ADC424B39FB6073D00D8048A31008017C1F826FFEF41FEEB027E3",
INIT_0B => X"7BEAF1C152201A4C05B7531D56B05B06A213FF863FF5D5F9FB5E8847A0702606",
INIT_0C => X"0D1030D1030D1030D1030D1030F0818688186B51BFDCC39732F3554866AD57C3",
INIT_0D => X"10080A20ED1D41880CC61A0044DFFC6EB5BCA06F18FC5A0E00F0038D1030D103",
INIT_0E => X"3FFE91FF98AEAA1AC6AC9A3A4AAD5B56ADAB56D5AFD572C597B147506203E8FC",
INIT_0F => X"0000260403C8948002000EC0000BC8948002000EC00010878AC3CB8AB8857202",
INIT_10 => X"EE0000400BC8948002000EC0000BC8948002000EC000097B0040200010003E02",
INIT_11 => X"400400003D80000070400DD81041400020003B80000410801AF0204180100000",
INIT_12 => X"010384008086378A080428C46A80080081002000780C800188000301017B0040",
INIT_13 => X"909042001C800409FC0020080001F80000007C0807484821000E400205D11101",
INIT_14 => X"10100A00003E020000BC0808EB01020280000F60000002BA222020407080102E",
INIT_15 => X"7520750000024080807868000100403C0808FA0040400000F8800001F02003F8",
INIT_16 => X"EF3AF6AF6389C2FE128971AB2DDDF8FFE0031B776BF4208006C0C92621F81000",
INIT_17 => X"D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B5",
INIT_18 => X"5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56",
INIT_19 => X"3FFFFFFFFFFFFFFFFFD5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D",
INIT_1A => X"0000001E0080397908000000A48710B4080240E543021B438A010825238B443A",
INIT_1B => X"4020100804020100800000000000000000000000000000000000000008200000",
INIT_1C => X"000A05028140A05028140A05028140A05028140A05028140A05028140A050080",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"8C2100804900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"02000100440408002408008002221000204116A280000F000001400000100010",
INIT_05 => X"00000000001265050080C000190002000000005C0000000A0000002C20600000",
INIT_06 => X"14016012000C405280200008001000011110012220009A88800009A880000000",
INIT_07 => X"0048912242288100800102000400010208000000040000082000002400814008",
INIT_08 => X"0A010040401080308400821155540001122448142491008A0049120408402210",
INIT_09 => X"04080A000000124058200408000880004440004080160C4100A8580099400000",
INIT_0A => X"4A50000080080E041000000008000C81000110010500002000000180001C8000",
INIT_0B => X"110091500020B408810000100200020408B0000020000081B2C208420ADA5353",
INIT_0C => X"5814058140581405814058140580A02C0A02C004800210C19808400500010009",
INIT_0D => X"10040860B188C0A80653020005A004039010280000800B00100040D814058140",
INIT_0E => X"600010000280000802050010660001000080004004900204020105302A000C42",
INIT_0F => X"0000A00000081480000001400000081480000001400000800C01082082210500",
INIT_10 => X"0000024000081480000001400000081480000001400000010000200000000000",
INIT_11 => X"4000000000000001400000080041400000000000000C00000010004180000000",
INIT_12 => X"0100000480802A40000000400000080081000000000000004800000000010000",
INIT_13 => X"1010420000002400040000080000000000024400000808210000001200010101",
INIT_14 => X"00100A0000000000028400004000020280000000000012002020204000009000",
INIT_15 => X"1000000000024080000000000010400400004000004000000000000510000040",
INIT_16 => X"8408420430E699AA42A1508104EA08000000810020000000044001AC20500000",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_19 => X"8000000000000000000010040100401004010040100401004010040100401004",
INIT_1A => X"20820800D41A8283AC618618EF1088160885001234B96061CCDEC4D205061170",
INIT_1B => X"6030180C06030180C08208208208208208208208208208208208208208208208",
INIT_1C => X"000B0582C160B0582C160B0582C160B0582C160B0582C160B0582C160B0580C0",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0803B2814D0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"26E1E905CC574828C4F85FC600000016004F77E2F887CDB80BC340DC07D1F000",
INIT_05 => X"F007E33E01D26CE43A92F2880B01F37011E93ED49BE01F1A03B8972E6D20F049",
INIT_06 => X"5AA06002026872BAE0B1282A005FFF001E1870223FC3BFC98101F109FC6780F1",
INIT_07 => X"3BC081023B233E804488527FDC008019968D74982C94110AF204001BC285A828",
INIT_08 => X"01E4191901A101B031F84000000831FA1028575A000110800124600C039C0020",
INIT_09 => X"C1111A0782082B50080508FF00048B124D4005C8AFF4154102914800110FFC00",
INIT_0A => X"B5AAF00A80A82C332D18ED301D229C82C7A93002017F405C409A42A9A51547F8",
INIT_0B => X"1158936D20601A98A10200308A002E240010BFC0600002AFFBE249420555A2A2",
INIT_0C => X"1A3401A3401A3401A3401A3401A9A00D1A00C000850400A11414C005005000B5",
INIT_0D => X"10080C60AB0F42A8046282000DBFFF13D059280201948B029029409A3401A340",
INIT_0E => X"6FFFF8000F8F80281A16A1504302058102C0816244B82A0CA25907D0AA015874",
INIT_0F => X"0080A40000283D80000001402000283D80000001402010901A7D694494192200",
INIT_10 => X"0000034000283D80000001402000283D80000001402002010000A00000000000",
INIT_11 => X"C000000000000081600002080341C00000000000008C00000410085380000000",
INIT_12 => X"81000006809076B2000040400001080581000000000000004810020002010000",
INIT_13 => X"1051620000003410040004080000000040026C00008828B10000001A00210909",
INIT_14 => X"00503A000000000042AC00044000228A8000000000801204212130400000D001",
INIT_15 => X"1000000001064180000000000010C02C000440000240000000000105B0001040",
INIT_16 => X"964C4A44A0C689FF3F9FFEC5D6DBFE0020096528A0B000000CC043EC60780008",
INIT_17 => X"6058160581605816058160581605816058160581605816058160581605816258",
INIT_18 => X"0581605816058160581605816058160581605816058160581605816058160581",
INIT_19 => X"17FFFFFFFFFFFFFFFFE058160581605816058160581605816058160581605816",
INIT_1A => X"AEBAEBFFF7FEFCFDF7FFFFFF5DE7CFCB773FFEFBFF3C7E1E779FFEFFF5060030",
INIT_1B => X"F7FBFDFEFF7FBFDFEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEB",
INIT_1C => X"000FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEF",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9E79E7BAF7DEBAFAFEFBEFBFFBFFDFFF7FCFF0FBFFDFF7EFDDFFFEFFE8000000",
INIT_1B => X"7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"0003F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"1084B030000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"6DA986092050306382C05A1C900000001FAE89016387B2A38B5000D03FA1C0C2",
INIT_05 => X"C0FFC338FF008048240426200081F147F1FB7F289B81FB8003A396D20940C3DB",
INIT_06 => X"098000C51000910100006C00426FFC7C202060445F1F2572060FE82671C607E1",
INIT_07 => X"0001020400440C41C000617FC0003021259CFDB01BF00020C001FF8040009800",
INIT_08 => X"2000200008020000000820440000100220489020000020000000000000000044",
INIT_09 => X"8004800E3CF3E0B1118C31747F000B33820209206FC9E80000000000220FD1FF",
INIT_0A => X"000687C0044040424B39FB6073C0010048A20000047C1F804FBEF01BEE8027E3",
INIT_0B => X"204A608142002A440492530C401049020221BF861FF0C06C493C800580000000",
INIT_0C => X"04003040030400304003040030600182001821011DCCC31222730048620C4382",
INIT_0D => X"000802004815010008840800405FF864008880661874500E00E0030400304003",
INIT_0E => X"1FFE81FF880EA000400098200C04080204010200810020C180904240400340B4",
INIT_0F => X"0000040403C0800002000E800003C0800002000E8000100780C2C30830806202",
INIT_10 => X"EE00000003C0800002000E800003C0800002000E8000017A0040000010003E02",
INIT_11 => X"000400003D80000020400DD01000000020003B80000000801AE0200000100000",
INIT_12 => X"000384000006118A080428846A80000000002000780C800180000201017A0040",
INIT_13 => X"808000001C800001F80020000001F8000000280807404000000E400001D01000",
INIT_14 => X"10000000003E020000280808AB01000000000F600000003A020000007080000E",
INIT_15 => X"652075000000000080786800010000280808BA0040000000F8800000A02003B8",
INIT_16 => X"223010010308025410082404A015F0FFE003182701B420800280C80201A81000",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_19 => X"17FFFFFFFFFFFFFFFFC080200802008020080200802008020080200802008020",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000080040",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"88280C4C7B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"00160090920C04800904848262220277E05152B280780D407428E723C01E1400",
INIT_05 => X"0F001CC000890026105810941C5C06800E008057641E00473C40680D32330C00",
INIT_06 => X"82541A028D584E40CB0583CCA0100000161F84322000DA8C40F003C80030780E",
INIT_07 => X"BF70E1C3BBBB1138AF7F888025340C0888430047040FEE182CA00044BC5827C5",
INIT_08 => X"CAFC1F1F07F0FE1C94F65B11555EAFFC1C306758B24197ABCDA467F2C9CF9B32",
INIT_09 => X"4FFB4730000011420A61080800B6E0C464258094101606D5A47A2A2098B02000",
INIT_0A => X"446000304A0488111084048E082D0ED020119D35F900002FB00105C01036D800",
INIT_0B => X"1FA599581D3A9583C105A892112C04C0A898403120071501A6C32222068A3050",
INIT_0C => X"789E07A9E0789E07A9E0789E070CF0184F038850A21008E514845AB510D0106D",
INIT_0D => X"9A95E954868AD0E52273F4AC2180000808061C01C48B0F81380CE0F89E07A9E0",
INIT_0E => X"4001120055704FC4A1624487E2489024481224091282C4300942A19439481842",
INIT_0F => X"5D65C3E3F01F52FFC1E0013C1F801F52FFC1E0013C1F8090423D38A18E3B15C9",
INIT_10 => X"118796BE001F567FC1E0013C1F801F567FC1E0013C1F9085DFBF7E15C06101C5",
INIT_11 => X"7E30F00C0270F3751F1FD00FECBF7E25C0700463E17B2C7F811FD7ADECC381C0",
INIT_12 => X"4190626D6491063597F9177B956EF378D33E4030061341F077C571F8F885DFBF",
INIT_13 => X"7F328E3082636B2807FFD80FE00007E03F7207D3E03F9167184131B5C40FE647",
INIT_14 => X"EFA0CAE06101C53E3647D3F144FCDD22B81C0098E57D9081FCE8C8520C4DAE20",
INIT_15 => X"1ADF08DBF81846A540049707E0FE3307D3F141FFB45478040570EED41F4FE047",
INIT_16 => X"C189601208A1502B4AA5584B4068000019A80098120BCA4C617635C938574FF3",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"A800000000000000000902409024090240902409024090240902409024090240",
INIT_1A => X"08208208831042720EE38E38AAF9C4C704DAB63A6D58B3C10BAE8E789AA09424",
INIT_1B => X"7C3E1F0F87C3E1F0F82082082082082082082082082082082082082082082082",
INIT_1C => X"0003E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F8",
INIT_1D => X"0000000000000000000000000000000030F007FFFFFFFFFFFFFFFFFFFFFFF900",
INIT_1E => X"155545F7AA975EFFFAABDE00FFAEBDFFF5D2EAAAAAF7AEBDEBA0000000000000",
INIT_1F => X"7FD5545FF8000155087FC0155F7D168B55007BFDF45085168ABA002E82145085",
INIT_20 => X"55568AAAFFFFD7545AA8028A00A2802AABAFF8028BEF5D7FFFE1000554214555",
INIT_21 => X"FFD168ABAF7AEAAAAAA2FFFDF4500043FE105D2E954BAF7FFC00100800175555",
INIT_22 => X"0002E974BA5D5168A00A2D142155005142010FFAE820AAFF842AABAA2AE95545",
INIT_23 => X"AAFF803FFFF5D2A821550000000BA007FD55FF5D7FC0145007FD740055041541",
INIT_24 => X"FFF082EBDF455D5142000082E82145FFD17DFEFFFD168BFFF780000BA007FE8A",
INIT_25 => X"FE3F000000000000000000000000000000000000000000000AAFBEAA00007BFD",
INIT_26 => X"6F0AA1C24AABEA495FC716F002A975FFE3AA95E00EBAEBDFD75D2AA8A80EA8E2",
INIT_27 => X"1FAE0016D56A16D557BC257D415E0216FA3F1E8FC0145B68B551475FAF6D1C55",
INIT_28 => X"7FEAA85487FD24AFE3D02DAAAE12BD5545A2803AA0000542A0070071C50BAFEF",
INIT_29 => X"B8A05A2AEA8B50F55A2F150005A3A438BD04AFAB8F550A8010E004924874825D",
INIT_2A => X"EA8A3AA05A2A5504001C74BA42A1571E8028E3DB7816D0120155EA568E870BAE",
INIT_2B => X"7ABA497A82FFAFD2A82485FD2415A105C21451ED42A002545E055FFBE81D0BE8",
INIT_2C => X"00B55EAAA100AA1D0F6F480B6A555A2A57A002A3D5FDB6A5C7E3DFFFE90B45B4",
INIT_2D => X"F45592E88A0AFE80A8B0A0000000000000000000000000000000000000000000",
INIT_2E => X"A1FD5D556ABEF5D557FEBA55022A3F70C6B405F4D2AE975EFAAAAB5E1AF3AABF",
INIT_2F => X"1CE0FDE69411A8DED57CE1055555E5F58EFFC01FE2CACB65F520EBE9EF67D7BE",
INIT_30 => X"034E0A592A4AD0079C75D6070CC5CBB0280C029ABAA3EBC11472800752117082",
INIT_31 => X"968BF57812A95E02A2AAB5EB0F280800EFAEE9F5D18F3142341D5DEEBEF55080",
INIT_32 => X"7D58AC448B69C30E02116220415A9540AA854140A0A2047F353AAF6C77F7F20D",
INIT_33 => X"56EEAB157ABEBE1B4D792A4AD1183454180DD3FDCAAAB7C91565455C141E4188",
INIT_34 => X"F0000001FF0000001FF01EABC4B8014174FF7DA80F52FEDE6BE93172D7D625B5",
INIT_35 => X"FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001FF0000001F",
INIT_36 => X"0000000000000000000000000000000000001FF0000001FF0000001FF0000001",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000100000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"CA1800080848B0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000010822C00803804000001999EF9C00040B0002000001000640200001018",
INIT_05 => X"08000000000100030008010468220A0004000000001000032000200002100800",
INIT_06 => X"8201961000060444010081002080000080820100000008004880000000284000",
INIT_07 => X"210C18306788C0089409800001140082000100010405000410A0000010082500",
INIT_08 => X"0A48903121780004C6000311555521F183060AC564BF818B5EDFDE0044600301",
INIT_09 => X"45B103200000140802234800000584000004808400020011A4581A2200002000",
INIT_0A => X"021000000800810400000402083000510000050020820036200005C00026C000",
INIT_0B => X"40000002000A008182200000002404400000000000010500008020A022220040",
INIT_0C => X"68064680646A0646A06468064690321503234204020018200404010784700404",
INIT_0D => X"C417C16004C0B838221090240180000801000C8800000190191064620646A064",
INIT_0E => X"6000000010200200802100022008100408020401020040100142200E0E08A20B",
INIT_0F => X"0021E300B000000781E00140018000000781E00140018000002430E30E0615C9",
INIT_10 => X"0000024E0000000781E00140018000000781E0014001908400005E11C0610000",
INIT_11 => X"3C30F00C000000155800D00000003E21C0700000000F00118000000468C381C0",
INIT_12 => X"40900004A400081401A0000004041218503E4030060000004804318008840000",
INIT_13 => X"01208C30800025200003D807E000000000725201600090461840001340002606",
INIT_14 => X"0F00C0E06100000012D2005100409520381C00000005920004C0C81200009A00",
INIT_15 => X"00120850B8180625400400000010711200510004B41478040000005548016000",
INIT_16 => X"40002002080000000804000A0000000011A000100208C008611430A000040250",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"0800000000000000000100401004010040100401004010040100401004010040",
INIT_1A => X"8A28A2AC8090C69606492492C09945235D5F7E2A5040B80E1C863A2958000500",
INIT_1B => X"DD6EB75BADD6EB75BAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A2",
INIT_1C => X"0002E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E975BA",
INIT_1D => X"00000000000000000000000000000000C0FFFFFFFFFFFFFFFFFFFFFFFFFFFC00",
INIT_1E => X"FE8BFF5D0002155557FFFFFF007FC21EFA2FFD74AAAAD5555550000000000000",
INIT_1F => X"D1574105D7FD75FFAAAA800AAF7AA974BAFFFBE8B45F7AEBDF455D2EAABEFF7F",
INIT_20 => X"5000015500557DF45AAD1400BAA2AE801550051555EFF7AA95400552AAAABAFF",
INIT_21 => X"F78028BFFFFFBEAB55F780020AAAA80020AA082EAAB5500517DF555D2EAAA105",
INIT_22 => X"5552A974AAF7AE820AA0851574BAA2D1574AA5D7BFDEBAFFD540155557FD5400",
INIT_23 => X"10557FFFFFFFFD56AAAAFFFFD7555AAD168B45AAAEAAABAFF842ABEF5D517DF5",
INIT_24 => X"E105D2E954BAF7AE80010082A97410557FEABFFAAFBE8BEFAAD1575EF557FFFE",
INIT_25 => X"056A0000000000000000000000000000000000000000000005D7FFDF4500043F",
INIT_26 => X"BDF55492AA8BC2EBDFEAF7F1F840017D4975D2FEF147FC51C7A2FBD5490BFD1C",
INIT_27 => X"4924385FAAA8AAAE3D145410F7F1D55D71C002DABAEBAA974BAF7FFEFB45FFAA",
INIT_28 => X"DB7DF7F540E2AE85028B40155145F7AF6DBED5450AA1C2080BEF495FC71D5412",
INIT_29 => X"FD56F16D5571D2E28E38E0216FA2D1E8E80140F45082B4002D082082AB8B6DBE",
INIT_2A => X"487BC70BFA97F7AF6D417E92482BF84020BA495557E3FF78E021FF1471FDEAAF",
INIT_2B => X"FF6FFD7FC7002FD74951D71EDFFABFD16FAAAE92BD5545A2DA3FB7DAAD4AAAAF",
INIT_2C => X"00547AB8F550A8010E00492487482FFFE82A85EBAE2FFC55554ADBD7A2FFC7BE",
INIT_2D => X"545AAFBF7400FBF9424F70000000000000000000000000000000000000000000",
INIT_2E => X"74AAF7FFFDF55F7AABFF55082CA8B4DF6C1E8F5E5400021EF005162BEF047FD5",
INIT_2F => X"225FF5843404547184164AA5D2EBEEB0A2D555410D3555714F8338AAAA1D0AE9",
INIT_30 => X"409000512AEABFFDF79DCBF755962010BDCBBC21455D7FEABEF75550ACBB7582",
INIT_31 => X"0688E5405D57D412F7D55F5E50C7F401BAAE8403CF5A3FFEAAEB083BC1000FF8",
INIT_32 => X"BD5FFE55F2AA9FEAFDF7F431A9F7FFE81FF013A8001AFF801F8BA0C57740BDAA",
INIT_33 => X"DA403FFFDA2FBF7FED2C7F955445079E280A00C56145EF5D16BABAA3EBC3157A",
INIT_34 => X"0000000000000000000596EBEF55080034E0A592A4AD00FB863550229BCABEB7",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000100000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0812",
INIT_01 => X"A145A00810790848048044A54E404340404000720885800802000906E4910200",
INIT_02 => X"5C010802020408040C455850AA055254090541A111200A104A0000000908B510",
INIT_03 => X"182002200C00004485264A001214912803150020218808002440854288890550",
INIT_04 => X"210302048014100160806B08702010102722C9E0412200651102418214049492",
INIT_05 => X"88510910540008812C06010018204342A58A08011290A1120A81230240018DCA",
INIT_06 => X"47450000022480090000210002A54C282122040CC9082D530085224410AA4204",
INIT_07 => X"2101020423408900940C402A900011012D41D518044C10025000AA8A50043D00",
INIT_08 => X"214912534123010085008010141521F020409260000100A00004428808102010",
INIT_09 => X"519D12041551589141A539C42A4C9608080004801700D10100311820A848E0AA",
INIT_0A => X"0244C28C000002025A81AE3048321002A700200900160AE42CAA839AA90442C1",
INIT_0B => X"42300225604004D080251121D0000400880178044355940A498C400004A00545",
INIT_0C => X"4F240472404F240472404D240441200692022B41365E53340EC6940564D012D6",
INIT_0D => X"00000620500403080A919000038AD03001C5080D1108C1009001404524045240",
INIT_0E => X"02AA40AA902408000010002220040C000201030201200C818098402082020438",
INIT_0F => X"0080A0000140000002000140200A8000000200014020100280E469C698353000",
INIT_10 => X"000003400A800000020001402009400000020001402008700000000010000000",
INIT_11 => X"0004000000000081400004C00000000020000000008C000010A0000000100000",
INIT_12 => X"0000000680004188000400840080000000002000000000004810000001420000",
INIT_13 => X"0000000000003409280000000000000040025000030000000000001A05100000",
INIT_14 => X"000000000000000042900000A100000000000000008012A2000000000000D026",
INIT_15 => X"4420300000000000000000000010C010000098000000000000000105400002A0",
INIT_16 => X"126000808200505448342228120090554000E00000000000088000A000000000",
INIT_17 => X"004010040300C0300C0300C0100401004010040300C0300C0300C01004010240",
INIT_18 => X"0400004000040000C0200C0200C0200400004000040300C0300C0300C0100401",
INIT_19 => X"9FC0FC0FC1F81F81F800C0200C0200C0200400004000040000C0200C0200C020",
INIT_1A => X"0410411823A4301040B2CB2CBACB002009C6B860185AA1491B0E2863E8001100",
INIT_1B => X"4A25128944A25128941041041041041041041041041041041041041041041041",
INIT_1C => X"03F25128944A25128944A25128944A25128944A25128944A25128944A2512894",
INIT_1D => X"00000000000000000000000000000000F0F007FFFFFFFFFFFFFFFFFFFFFFFC07",
INIT_1E => X"415410AA8415555087BFFF55A2AA800BAFFAE9540008002AA000000000000000",
INIT_1F => X"FBEAABA5D7FE8B555551421455D0002145552EBFEBA007FC21EFA2FFD75EFAA8",
INIT_20 => X"2AA974BAFFFFE8B45552EBDF45FFAEAABFFF7FFE8B55F784155EFA2AEBDEAAA2",
INIT_21 => X"5D7FFFF555D2AAAAAA5D2E820BAA2FBEAB5555557DF55A2AEBDF555D2E954BAA",
INIT_22 => X"55D043DEAA5D04021EF557FC21FFAA8428BFFAAAA954AAAAAAAAAAAFFD157410",
INIT_23 => X"FFA2D17DFEFF7800215500557DF55AA80001FFAA80001550055575EFFF840215",
INIT_24 => X"0AA082EAAB5500517DF555D042AA10A284154005D0015410085568A00FF80175",
INIT_25 => X"8A2A0000000000000000000000000000000000000000000005D00020AAAA8002",
INIT_26 => X"C51C7A2FBD55D2BE800042AFE8E1557D0075D2F45BEAA800AAFFAA9543A08003",
INIT_27 => X"0105FFBC20BDEAAA2FBF8AAA557BE8B6D5D5FFABEF49040017D5D20B8EAA007F",
INIT_28 => X"A0BDF7D480E174BFA02A974BAF7F5EFB455D2ABDF55492AA8BC7EBDFEAFEFFD0",
INIT_29 => X"6AAADAAAE3D155E105571D55D71C002DABA5524820BAB6FFEFB6D555578F7DB6",
INIT_2A => X"0155C51D0092A071555D5E3AE821D00001FF0871C016DBED1FDE90E3A497492B",
INIT_2B => X"8007FED000E3DA3DFD5E3DFFFBD5A38A021551C5F7AF6DBE8F401D7B6A000147",
INIT_2C => X"00410F45082B4002D082082AB8B6D1C5B7DF7FF78E075C5BE8555400550A3842",
INIT_2D => X"0AAF7AA954AA00042AAA20000000000000000000000000000000000000000000",
INIT_2E => X"21EF55042AAAA007FD5555AAFBD7545FBB8020A3F7AE975EF005560B55F7AA80",
INIT_2F => X"A8F45A6C1E8F5EFF84165EFF7802BAB0A2FFEAABA557BEABEF057D68F5F5A000",
INIT_30 => X"BFFFEF04552ABFFFF841FFE75CA882108202E974AAF7D57DF55D7AABFF5428AC",
INIT_31 => X"D1E00A1A884174A8FFAEBFEB0A2D55541051555694F002CA8AA80800020AAF7F",
INIT_32 => X"680800FFF7AAA155F595542455512A975455D3AA8A005500151FF0C57401E5F3",
INIT_33 => X"7895554005D2A8A0B882FFFFE10AAAAAB755A66B6AF56A2AA801455D7FE8BFFF",
INIT_34 => X"00000000000000000000C3BC1000FF8409000512AEABFF5D79FCAF774AE005BE",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000200000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380206",
INIT_01 => X"014C9A40408001683C0462C99E004B61404040028804A0080A000D16A0990A0C",
INIT_02 => X"4809A902031800444460589C66E331352180D468B8240E600C0081110B80ACD0",
INIT_03 => X"DA14C2210C0001D235834A0648D60528330006810A80881068A80C029CC56330",
INIT_04 => X"20886819A02740ECD2107364B37569100A04C1E01CA52010990240420E205A08",
INIT_05 => X"5831803532410000260E272058232259954369000A506912018CA582480038D1",
INIT_06 => X"8381A014000200AC2190ED0002ACD99881822144C5A409430682800046294140",
INIT_07 => X"218408142740E2C0948C3066500071913209CC8004640102D003999552083D20",
INIT_08 => X"00409231296AA180C2000110001521F0810A92E7402F00AB0016CA080C600111",
INIT_09 => X"41B112014D30E43802A76DD09905882B010605A01A4941010211088A2A43A399",
INIT_0A => X"4A12D9820880832264119D004860900104002008000F399606BC07998BA546AC",
INIT_0B => X"42522013604080D084A01001C8302D00008153000731C3000988C0040A224110",
INIT_0C => X"602406824068240602406224068920151203030032545B7404D7804566594796",
INIT_0D => X"080600E04C442068088590000999C8E84041086C001091009001406824060240",
INIT_0E => X"E6660599902600209021204A010E1C850C428521C208480021D842081A03E231",
INIT_0F => X"0090000003200000000010002008A00000000010002008038666928B28A65300",
INIT_10 => X"000801000A200000000010002009E0000000001000200A380000000000000000",
INIT_11 => X"0000000000000088000002D00000000000000000028010001620000000000000",
INIT_12 => X"0000008201021C88000048800280000000000000000004000010000003600000",
INIT_13 => X"8000000000041019980000000000000040802000068000000000020805B00000",
INIT_14 => X"0000000000000000C020000C8300000000000000008200AE000000000010402B",
INIT_15 => X"41003100000000000000000002008020000C3800000000000000012080001298",
INIT_16 => X"737420C20A01405468360022201185CCE0128410820000008088021C40A00008",
INIT_17 => X"2108721085218852188521885218852188521887210872108721087210872308",
INIT_18 => X"1086214872108621C852188421C852188421C852188721087210872108721087",
INIT_19 => X"26AA555AAB554AAB5561C852188421C852188421C85218842148721086214872",
INIT_1A => X"0410412881D0B0000092492480A981E063C638321450A08899A62C314A810508",
INIT_1B => X"EA753A9D4EA753A9D49249249249249249249249249249249249249241041041",
INIT_1C => X"BC4351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A9D4",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF82A",
INIT_1E => X"02AA00AA843DF55FFAA955EFA2D168B55557BEAA000055420000000000000000",
INIT_1F => X"5568A00087BE8BFFA2D155410AA8415555087BFFF55A2AA800BAFFAE95545080",
INIT_20 => X"D0002145552ABFEBA007FC21EF007FD75FFAA841541008002AB55AAAA955EF00",
INIT_21 => X"5D7FC0155005168B455D042AB45F7FFD741000042AA10AAAABFF5508003FF555",
INIT_22 => X"A5D7FC2010A2D1575FFF7AA975555D2E80145F78415545082EBDEAAA2FBEAABA",
INIT_23 => X"FFFFAAAAB55552A954BAFFFFE8B55552EBDE00F7AEAABFFF7FBEAB55F7AABDEB",
INIT_24 => X"B5555557DF55A2AEBDF555D2E954BA002EAAABA002A821EF5555554AA087BC01",
INIT_25 => X"203A000000000000000000000000000000000000000000000082E820BAA2FBEA",
INIT_26 => X"800AAFFAA95578080038A2AA28E3AF55E3A0BA5D7AADB6FB7D5D7FEAA3808554",
INIT_27 => X"E2AB55B6A0925D7085F6AA10087FEABD7AAD57AEBAB68E1557D1475FAF45BEAA",
INIT_28 => X"AEBFF6D1D04AAFFA41040017D5D20B8EAA007FC51C7A2FBD55D7BE80004AA1E8",
INIT_29 => X"C20B8EAAA2FBE80AA557BE8B6D5D5FFABEF49002FB55FFF5D0438140E2FA38B6",
INIT_2A => X"EBDFEAFEFAB8ABAE925D21C7010EADB525D7FFAE975C75D0A901FFFF801557D1",
INIT_2B => X"74971D24820875C21D5EB8AA8FFF012A954BAFFF5EFB455D20BDE00EBAAA8BC7",
INIT_2C => X"001C24820BAB6FFEFB6D555578F7DB6A0BDF7DEB8E125FF002EADA921420871D",
INIT_2D => X"FFF5D7FEAABA0051400A20000000000000000000000000000000000000000000",
INIT_2E => X"75EF555168B55F7AA800BAF7AA955EF00042AAA2A2AEAAB55A28408145AAFFFF",
INIT_2F => X"D7145FBB8020A35D2ABEF55F7800015F087FEAA00007FEAB55FAD568AA2AFAE9",
INIT_30 => X"5420BA5D2ABFEAAF7AE9DFF759A82AEF70800021EF55042AAAA007FD55558A7B",
INIT_31 => X"040255FFD84175EF55002AAB0A2FFEAABA557BEA3EF057968F575D003FF55F7D",
INIT_32 => X"52A3FF10AA8429F45A7D5EAF5FFBAEAAA10554155400AAFFD5145FBAC9755F05",
INIT_33 => X"052ABFE10550415557085540000005156155FE90A8F5C082E974AAF7D57DF455",
INIT_34 => X"00000000000000000005500020AAF7FBFFFEF04552ABFFFF843FFE77C80825BC",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000100000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10804002061080A284201081034809800A00230340007833522C82D04A16002",
INIT_01 => X"80439982183828490400050E12000340403008418984014902030106A0D10204",
INIT_02 => X"480108A000000000446418E01E80F00A41043118680402000800000009882390",
INIT_03 => X"0CA080210C0000408006480002001120260012603000000030808900888100F0",
INIT_04 => X"4403A609A055306B82C0705800CEE510082AC0A16B0350E3808041D03865D002",
INIT_05 => X"C0F20B36F0000901240626200820E26780E244A19A41E4020BAB06404001D312",
INIT_06 => X"434420151220118900806922406C3C7800201448DD9D2870020F228075A60715",
INIT_07 => X"2181000023480040840C001E180030032009700024641002C00187A440047C00",
INIT_08 => X"084830110160208004000001101121F220000260000100AA0004408000000001",
INIT_09 => X"519102063DF3E02B100B097407448F200A0209A041CA290102130C8800466478",
INIT_0A => X"8543D048006040064010E4007F62110105002002044007846124E0A00E0DC1EB",
INIT_0B => X"60020291404024808030512C40106D022203B1445810856A019400058F8404B5",
INIT_0C => X"052430D24305243052430D24304121A6921863013FD8807626EE000D64540284",
INIT_0D => X"28081080508104400A00800009B878680000880C1160410C90C143152430D243",
INIT_0E => X"81E0E18790012A00080102280800000202010102810020018098404110020004",
INIT_0F => X"0090000005E0200000001000200C6020000000100020000390E6C30830806204",
INIT_10 => X"000801000D20200000001000200EE0200000001000200A6A2000800000000000",
INIT_11 => X"8000000000000088000003B00100000000000000028000002EA0001000000000",
INIT_12 => X"80000082000251D80000C0044280000100000000000004000010000003282000",
INIT_13 => X"00002000000410121800040000000000408030000B8000100000020806F00000",
INIT_14 => X"0000100000000000C030000C9000008000000000008200FC000010000010403B",
INIT_15 => X"A500100000000100000000000200803000042E000200000000000120C0001590",
INIT_16 => X"30000800002400044934040AA231B63C20530801000410009889821040A00008",
INIT_17 => X"00401008000040300800004010000200C01000020040100802004030000002C0",
INIT_18 => X"000000C0300401008000000200C0100C01000020080000C030000000C0100802",
INIT_19 => X"325930C9A6CB261934C000200800004030040300800000020040100C03000000",
INIT_1A => X"8A28A2BD30264686668A28A2605145031C03F028000A1C2ED7831A2820244140",
INIT_1B => X"8D46A351A8D46A351AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA28A28A2",
INIT_1C => X"CFB068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D068351A",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF82B",
INIT_1E => X"54200000557FE10FFFBEAA10007FD7410FFAA97555082A800AA0000000000000",
INIT_1F => X"043FEBA5D7FEAA00007BE8AAAAA843DF55FFAA955EFA2D168B55557BEAB45005",
INIT_20 => X"A8415555087BFFF55A2AA800BAFFAE9555508002AA000055574105D2A800AA00",
INIT_21 => X"087BE8BFFA2D17DE1000517FE10AAAAA8AAA002E97545557BC00AAA2FFEAAAAA",
INIT_22 => X"0F7FBC2010A2D157400AAAE974AAAAAA974BA08002AB55A2AA955EF005568A00",
INIT_23 => X"AAA2FBD54BA080002145552ABFEAA007FC21EF007FD75FFAA8417410A2D14000",
INIT_24 => X"41000042AA10AAAABFF5508003FF55F7D568A00552EA8BEFA2AABDEAA087BEAA",
INIT_25 => X"50B800000000000000000000000000000000000000000000055042AB45F7FFD7",
INIT_26 => X"6FB7D5D7FEAB7808554203A145178E00FFFBE8A101475D5400F7A49057D08248",
INIT_27 => X"157428492E8008200043FE925571EFA380871C7028A28E3AF55F7A0925D7AADB",
INIT_28 => X"75C5092AAF5FDA38BE8E1557D1475FAF45BEAA800AAFFAA9557D080038AAA145",
INIT_29 => X"6A0925D7085F6AA10087FEABD7AAD57AEBA08517DE00AAAEA8A9200249056D41",
INIT_2A => X"BE80004AAFEDB42028EBFBC2028BED152438AAA092492AAA4954281C0E2FB55B",
INIT_2B => X"FAA803DEBA0875EDA80BEF1C743840040017D5520B8EAA007FC51C7007BD55D7",
INIT_2C => X"0041002FB55FFF5D0438140E2FA38B6AEBFF6DBE84AAEBAF7DF6AA00412EAABF",
INIT_2D => X"410FF84021EF0800154B20000000000000000000000000000000000000000000",
INIT_2E => X"AB55F78400145AAFFFFFEF5D7FEABFF0051400A25D5568A00FFFFEAA105D5155",
INIT_2F => X"955EF00042AAA25555410BA082E8201000043FE005D517DEBA0851574B2AAAEA",
INIT_30 => X"AAAA000804001FF005575408AA557FEB2FFAE975EF555168B55F7AA800BAF7AA",
INIT_31 => X"AC154B25F2ABFF55F7800015F087FEAA00007FEAB55FAD568AA200557DE00AAA",
INIT_32 => X"07FD5555087BD6145FAAC000A2A6FBC00BAAAFBC00BAF7D1550AAAA8002010F2",
INIT_33 => X"F7FBE8A00082EA8BFFAA843FEBA08517DE00F3F9574B30800021EF55042AAAA0",
INIT_34 => X"000000000000000000008003FF55F7D5420BA5D2ABFEAAF7AEBDFF779A82AA43",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000200000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF0A0791B3FC1694378283C81FD996A091A32142007A336A20E03C040C002",
INIT_01 => X"A91FBDC4983088485C4A60000C24C26041280A00084000C8C212812EE2953231",
INIT_02 => X"C809AD5EB118E640A4F548FC011FF0002080000082ECC66609DB7DDDCB1FA036",
INIT_03 => X"4A120E4D3E4C90D294A31E824A52847A0B20640A88800000B8E0FD522885500E",
INIT_04 => X"001440849A2604001934800041110A71E2B068B110DB321C662AE22DC08A3448",
INIT_05 => X"370C14CA0E0800022446011C4E7F17907BEBD1AA65AE10571450DFC152522449",
INIT_06 => X"07319A109D129D450A846FE4E24C0305A1A5901C82416D05417118630839B88A",
INIT_07 => X"A5B56AD5A718C038AFFEA9FE39348C9204C389672407EE120EA5806E6C503AC5",
INIT_08 => X"C05896372728FF8C420619000003AFF4AD52A2C5D26F0EABCC96CD7AC4639902",
INIT_09 => X"5BD3571182080C000041080300F6F0C72221889C6FE20395A013282002B029F8",
INIT_0A => X"A23D203042444124098516CE0C2D13512410AD3CF8014005902DA6B2D1A4D810",
INIT_0B => X"645528937D5A85D3C4B0F883C10C24E0022B0E310612C2684CA16320A60A1185",
INIT_0C => X"288E3388E3208E3388E3288E330471904719C31438D04930ACE40FFD727C4304",
INIT_0D => X"8297A454544032252811E4AC2387F91008839C6CC413958D38C4E3208E3308E3",
INIT_0E => X"7FE0627FC25847C421516685844480204211200810028C38089AE00C894AA201",
INIT_0F => X"5D65E1E3C037E37FC3E0017C1F8037E37FC3E0017C1F900040261083080610CA",
INIT_10 => X"118796FE0037EA7FC3E0017C1F8037EA7FC3E0017C1F9300DFFFDE15D06101C5",
INIT_11 => X"BE34F00C0270F3754F1F8207FDBEBE25E0700463E17F3C7E054FF7BE6CD381C0",
INIT_12 => X"C090626DE40150459759573BBD6EF37D523E6030061341F07FC570F8FA00DFFF",
INIT_13 => X"6FE2AC3082636F301BFFFC07E00007E03F7263D383B7D1D6184131B7C1FEF64E",
INIT_14 => X"FFA0F0E06101C53E36E3D3EC84FDDDA8381C0098E57D923FDFC8D8120C4DBE0B",
INIT_15 => X"6FDF58DBF81C072540049707E0FE7323D3E43BFFF61478040570EED58F4F9397",
INIT_16 => X"00C108901822490448260224000040FC390250A2110B8ACC48B206A159A74FAB",
INIT_17 => X"08422080210882108C220842008821088230842208C20088210802308C2008C2",
INIT_18 => X"8422080230882108823080230842008C22084220842008C20080230802108C20",
INIT_19 => X"1092596D34924B2DA6884220842008821080230802108821084220842208C200",
INIT_1A => X"BEFBEFB7F7FE7EFEEE79E79EFAF2DDA73FBDCEDBFF9D3F0FDE0DB6DBF4208506",
INIT_1B => X"F77BBDDEEF77BBDDEEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"FED7BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF804",
INIT_1E => X"A800AAAAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF0000000000000",
INIT_1F => X"7FD7555A2D5575EF55517FF5500557FE10FFFBEAA10007FD7410FFAA97410082",
INIT_20 => X"A843DF55FFAA955EFA2D168B55557BEAB55005542000007FD74000055574BA5D",
INIT_21 => X"5D7FEAA00007BC00AAAAAEBDF45A28428B45FFD168BFF00002AABA5D2ABFFFFA",
INIT_22 => X"0F7D57FEBAFF80174BAAAD1555EF5555555550055574105D2A800AA00043FEBA",
INIT_23 => X"BA557BD75FFAA8415555087BFFF55A2AA800BAFFAE95555080028A00A2FFFDE0",
INIT_24 => X"AAA002E97545557BC00AAA2FFEAAAA082A97545F7D5420BA5D2E821FFA2D5554",
INIT_25 => X"DFEF00000000000000000000000000000000000000000000000517FE10AAAAA8",
INIT_26 => X"D5400F7A49043D0824850B8A2AE9756D145B401FFFFFFC7010BEDF524AA5571F",
INIT_27 => X"1D74380851524BA5571D757DB6D5525EF555178F6D145178E00EBFBE8A101475",
INIT_28 => X"0A28AAA5524BFFFFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D0855420BA147",
INIT_29 => X"92E8008200043FE925571EFA380871C7028B6AEBDF45B68A28B6DEBDF6DBEF1C",
INIT_2A => X"080038AAAA2FBF8E10EBD578EAAFF8415482BED1555EF55555057D1451524284",
INIT_2B => X"A552A821FFB6DF574A85575C55EFBE8E1557D1475FAF45BEAA800AAFFAA9557D",
INIT_2C => X"0008517DE00AAAEA8A9200249056D4175C50920875FDA381C209256DFFDF420B",
INIT_2D => X"400F7FBC00BA55557DFF70000000000000000000000000000000000000000000",
INIT_2E => X"8A00AAFFEAA105D5155410FF84020AA0800154B2AAAA975FF5D7BC21EFF7FBD7",
INIT_2F => X"EABFF0051400A25551554BA0051400BA5551575EFF7D1401FF5D5568BE755556",
INIT_30 => X"AAABFFAAFFFDFFF552EA8AAA55043DFF7AAAEAAB55F78400145AAFFFFFEF5D7F",
INIT_31 => X"55421E75555400BA082E8201000043FE005D517DEBA0851574B2FFAABFF45FFA",
INIT_32 => X"7AA800BAF7AA955EF00002AAA2A2FBE8A00A2D16AAAAFF8002410FFD5575EF55",
INIT_33 => X"5D00021FFFFFFC00BA552A821EFFFFFD74BA5D51575F7FFAE975EF555168B55F",
INIT_34 => X"000000000000000000000557DE00AAAAAAA000804001FF0055554088A557FEB2",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000C00000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C03002818000400322120040B313301C4389B2082",
INIT_01 => X"A74041CA38396849188160000C42424041000000090800090210090008110200",
INIT_02 => X"080108200C1000004465580000C0080100000000010432400800800009882050",
INIT_03 => X"080200010C234040842248600210812183806504488000103080014E88810000",
INIT_04 => X"0040504288A68210003120000000001002A0E8A910A072101000400A00203040",
INIT_05 => X"2800000400241801A52500094A02022014100128005004020010A1C044C02800",
INIT_06 => X"232000044084804914CA7C011AA3FC012122104CC0812D403280182308294000",
INIT_07 => X"2181020423488002940C0401D0480112000100004404004602447F8051223912",
INIT_08 => X"004812130160008304000000000021F020408264000108A00004400030400000",
INIT_09 => X"419102010104000A100348037F0584230A902A894008090343108802000FF407",
INIT_0A => X"B22D77C12052522400000400883011210000220006FC5FA400401484002447E0",
INIT_0B => X"60422291504420D084B0502044811428222300004611C57849A0150CA98A8561",
INIT_0C => X"1025B1025B0825B0825B1825B1112D8012D803003AD0413424E4014D627C0704",
INIT_0D => X"4404074040900B300A00810001A0021825E0886C0110916C96D15B0025B0025B",
INIT_0E => X"001E0800122100120499210A04A54652A12850962945180A14B44002CC020080",
INIT_0F => X"008ABA0030202100000001402068202100000001402067401026000000000031",
INIT_10 => X"00000341E8202800000001402068202800000001402062840000800000000000",
INIT_11 => X"8000000000000083D00052000100800000000000008CD0018400001200000000",
INIT_12 => X"800000069A48584000A0400000000005000000000000000048128D0002840000",
INIT_13 => X"80402000000034C1E000040000000000400FE000644000900000001A34000008",
INIT_14 => X"00003000000000004BA000112B0000880000000000807E80010010000000D1A4",
INIT_15 => X"0020250000040100000000000010CCE000198000020000000000010F80006028",
INIT_16 => X"0A728CA8C22540444924050CA9120603E0A2024048400010298432A002A00050",
INIT_17 => X"94E519465094A53946519425094A53946509425294E53946509425394E539625",
INIT_18 => X"425294E509425194E5294A519425094E5394A509465194A5294A519465094A52",
INIT_19 => X"3B1C618E38E38C31C71425294E53942519465294A53946509465394A50946519",
INIT_1A => X"8E38E39DB3B676F66EFBEFBEFAFBC5E73FC7F87A7D4ABFE7CFAFBE7BFA05004A",
INIT_1B => X"7F3F9FCFE7F3F9FCFE38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E3",
INIT_1C => X"6B23F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"00000000000000000000000000000000C0F007FFFFFFFFFFFFFFFFFFFFFFFC08",
INIT_1E => X"FFDFFF087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF0000000000000",
INIT_1F => X"AA97555A2FBD7410AA8428AAAAAAE955450055421FFFFFBC0010AAD5574BA557",
INIT_20 => X"0557FE10FFFBEAA10007FD7410FFAA97400082A800AA08515555508043FE00F7",
INIT_21 => X"A2D5575EF55517FF55A2AA97400552AAAB45082E80155F7D1575EFFFAA955550",
INIT_22 => X"0FFD5401FFF7AAA8A10082EAAB45A2FFC2000007FD74000055574BA5D7FD7555",
INIT_23 => X"BAFF843FFFFAA843DF55FFAA955EFA2D168B55557BEAB5500554200000003DE1",
INIT_24 => X"B45FFD168BFF00002AABA5D2ABFFFF087BD5545007BFDE10AA803FE105D516AA",
INIT_25 => X"25FF000000000000000000000000000000000000000000000AAAEBDF45A28428",
INIT_26 => X"C7010BEDF524AA5571FDFEF1C7BFFF55FFA095482B6A49256DEB84104BAFFD15",
INIT_27 => X"B5057D1C003DE28F7A49057DAAF5D2428A2842AAAAA2AE9756D145B401FFFFFF",
INIT_28 => X"DF525FFFFA49756D145178E00EBFBE8A101475D5400F7A4904380824850381C5",
INIT_29 => X"851524BA5571D757DB6D5525EF555178F6DAAA495428412AAFB451C2A8017DE3",
INIT_2A => X"0855420BA1C0E3FE00E3DB471EFE3AAAAA00082EA8B6DA2F1C50381471D74380",
INIT_2B => X"0A28038E1049516AAB8FF8428FEFA28E3AF55F7A0925D7AADB6FB7D5D7FEAB7D",
INIT_2C => X"00B6AEBDF45B68A28B6DEBDF6DBEF1C0A28AAA5524BFFFF1C7BD057D1C71FFE1",
INIT_2D => X"1FFAA84000AAFFD1401E70000000000000000000000000000000000000000000",
INIT_2E => X"75FF5D7BC21EFF7FBD7400F7FBC00BA55557DFF7557BFDF55F78017400F78000",
INIT_2F => X"020AA0800154B2557FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2AAAA9",
INIT_30 => X"ABDF555D2A821EFAAFBC01FFF780155F7555568A00AAFFEAA105D5155410FF84",
INIT_31 => X"D5554B25551554BA0051400BA5551575EFF7D1401FF5D5568BE7AA80174AA082",
INIT_32 => X"AFFFFFEF5D7FEABFF0051400A25D2EBFE10AAFFD55EFA2AEA8A10082EA8BEFAA",
INIT_33 => X"557BC01EF55557DE00AA842AA0000516AABAFF8428BE7AAAEAAB55F78400145A",
INIT_34 => X"0000000000000000000FFAABFF45FFAAAABFFAAFFFDFFF552EA8AAA55043DFF7",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000900000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0048201002842002C024500188000003000000003302300C018180006",
INIT_01 => X"020008402008404C042080000211024840000000080000080200010008110200",
INIT_02 => X"4801082248100000444008000080000041000000002222400800000009008010",
INIT_03 => X"0802010288A1484000020A400000002902006480088000003080040408810000",
INIT_04 => X"00004804890640004032030010000010008060E4100000140004500800403040",
INIT_05 => X"20000004004208016606010A0A20022000000000004000228010010080882000",
INIT_06 => X"030060004084004820906D311080020101000000008008011000000308290010",
INIT_07 => X"2100000023008002940C04000A4A010200018920646C10C50350002442003820",
INIT_08 => X"084812130160214204000000000121F000000244000100AA0004400920400000",
INIT_09 => X"419122810000081A00876882000590081100448A1000002350100CAA20002800",
INIT_0A => X"050280020100020400011640CC72602900044280028180242008069081244010",
INIT_0B => X"00200411508500B08805054C18024432A002400C99E410000080451100070014",
INIT_0C => X"05448054481544815448154481C22406A2406851201000200484950500F0145E",
INIT_0D => X"0144414A40000022880081511180036040044A013268E1205202480544805448",
INIT_0E => X"6000600010000020001102080102048102408120402800086098480008A20000",
INIT_0F => X"A2081210380021000001E003C0580021000001E003C042283426000000000021",
INIT_10 => X"00706801980028000001E003C0580028000001E003C044840000800009864038",
INIT_11 => X"80000330C00F0C0210807000010080000581C01C1C009201C000001200001607",
INIT_12 => X"8C2419101028D00020A2000000000005080082C180603A0E002A090404840000",
INIT_13 => X"8040204321188095F8000400061E001F800C202077C0009021908C4029F00008",
INIT_14 => X"00003009864038C10820201FAB000088026130071A00613E010011848322014F",
INIT_15 => X"6520350000640912058100F81C0108A0201FBA0002008239020F100880807BB8",
INIT_16 => X"114400C0002140144C2480200000040024A28400800044222980300CC4A0805C",
INIT_17 => X"2048120483204802008020082200812048120481200802008020081204812048",
INIT_18 => X"0880204812048020080200812048120080200802048320481204802008220080",
INIT_19 => X"2C208200010410400020C81200802008120C81204802008020C8120481200802",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000002A1050A",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"9840000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF818",
INIT_1E => X"5555FFF780155EFAAAEA8ABAAAFBFDE0055556AA005D04155550000000000000",
INIT_1F => X"AAAAB455D556AA00FFAE95555087BFDF45F7AA974AAAAAA97555F784174BAF7D",
INIT_20 => X"AAE955450055421FFFFFBC0010AAD5574BA557FFDFFF5555555EFAAFFFDFEFAA",
INIT_21 => X"A2FBD7410AA8428AAA557BFDFFF55003DFFFF7FBEAA00002EAAAAA082EA8A00A",
INIT_22 => X"FA28000010552EBDE00007BEAAAAA2D14000008515555508043FE00F7AA97555",
INIT_23 => X"55557BD55FF00557FE10FFFBEAA10007FD7410FFAA97400082A800AAF7AE975F",
INIT_24 => X"B45082E80155F7D1575EFFFAA955555D51574AAAAFFD5545087FEAB455D516AB",
INIT_25 => X"7555000000000000000000000000000000000000000000000A2AA97400552AAA",
INIT_26 => X"9256DEB84104BAFFD1525FFFF8E175C7A2AAAAA82A2F1FAE105D556AA10410E1",
INIT_27 => X"B575D7AAF1FFFD7AAAAAFB7D495F6AA10E3AE905551C7BFFF55FFA095482B6A4",
INIT_28 => X"2EA8A821C2EAAA00A2AE9756D145B401FFFFFFC7010BEDF524AA5571FDFEF415",
INIT_29 => X"C003DE28F7A49057DAAF5D2428A2842AAAA497BFAFFF49003AFEFEBFBEAA001C",
INIT_2A => X"082485038F7A4905C7A28A070384120BDE100075EAA82BEDB470101C5B5057D1",
INIT_2B => X"5087BE8B7D555F6AB57417BC05D7145178E00EBFBE8A101475D5400F7A490438",
INIT_2C => X"00AAA495428412AAFB451C2A8017DE3DF525FFFFA49756D495150492BEF1D255",
INIT_2D => X"A00555168A10002E9754D0000000000000000000000000000000000000000000",
INIT_2E => X"DF55F78017400F780001FFAA84000AAFFD1401E7FFAA97555A2AEA8A10AAD568",
INIT_2F => X"C00BA55557DFF7007BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215D557BF",
INIT_30 => X"028BFFAAFFEAA105D2EAAA005D2AAAA18AAAA975FF5D7BC21EFF7FBD7400F7FB",
INIT_31 => X"FBD7408557FC01EF55043FEAAFF80021EFA2D1420BAAA8428AA2007FE8BFF080",
INIT_32 => X"D5155410FF84020AA0800154B2FF8402145A2AA954AA00043DE0000516AA10F7",
INIT_33 => X"005140000FFD140145007FE8BEF557BEAB55087FC215D555568A00AAFFEAA105",
INIT_34 => X"0000000000000000000AA80174AA082ABDF555D2A821EFAAFBC01FFF780155F7",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"A140084000080048040100000202024040000000180800080200010048110204",
INIT_02 => X"080108020090000004655C000080000051000000002402400800000009008010",
INIT_03 => X"0002000100300C408422420002108108028065844880001030808D4288810000",
INIT_04 => X"0002584288A2C210003103001000001002A0E8C910A032541000090A00643040",
INIT_05 => X"2800080400645049A725010942220020140001A9005000004810A0C0044D2800",
INIT_06 => X"630400041404B141345A7C00426FFC01292214444081254102801A2308214004",
INIT_07 => X"21810204214080069408000008C3010200018920E06C0000021DFFA453263D32",
INIT_08 => X"084010110120018024000000000021F020408264000000080004400802400000",
INIT_09 => X"51B1004100040898128768820045142B0B902E895008080A1B13848A20002800",
INIT_0A => X"522920032052520400011641C460010D000000C8040100260008061081204010",
INIT_0B => X"4262229150012080102500211C81142880224000400411784920410C208514A4",
INIT_0C => X"0020000200002000020000200011000810008A55201000200484950004F0145E",
INIT_0D => X"40284301481509004885900101A0020964240109011890008011001020000200",
INIT_0E => X"0000200002210A320489000005A142D0A16850B6294D100A34B05242401340B4",
INIT_0F => X"00800008100001003C1FE00020080001003C1FE0002004401424008208041001",
INIT_10 => X"00000100080008003C1FE00020080008003C1FE000200080000001EA2F9EC000",
INIT_11 => X"01CB0FF3C000008000201000000081DA1F8FC0000080110080000002132C7E3F",
INIT_12 => X"3E6C00020040480040200000001004862CC19FCF81E000000010000200800000",
INIT_13 => X"004C11CF60001018000003F01FFE00004000000420800688E7B00008042000B8",
INIT_14 => X"000F251F9EC00000400004050002005D47E3F00000800084011607AD80004021",
INIT_15 => X"0000822406E5B85A3F830000000080000405000009AB87FB0000010000103000",
INIT_16 => X"1A768C68D260001448242704B912040002200640484000110104300042002018",
INIT_17 => X"B46D1B46D1B46D1B46D1B46D1B46D0B42D0B42D0B42D0B42D0B42D1B46D1B66D",
INIT_18 => X"46D1B42D0B42D0B42D0B42D1B46D1B46D1B46D1B42D0B42D0B42D0B42D0B42D0",
INIT_19 => X"200000000000000000346D1B46D1B46D0B42D0B42D0B42D0B46D1B46D1B46D1B",
INIT_1A => X"9E79E7B7F11E66C6FAD96D96520145052A1F5E2BD085122ED48F3AEB20840442",
INIT_1B => X"1F0F87C3E1F0F87C3E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"A6D4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87C3E",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF805",
INIT_1E => X"415555080000000087BEAA10F7803DE00FFAEBFFFF0800155FF0000000000000",
INIT_1F => X"80154105D7FC2145005155555F780155EFAAAEA8ABAAAFBFDE0055556AA005D0",
INIT_20 => X"87BFDF45F7AA974AAAAAA97555F784174BAF7D5555FF552AA8AAA557FC0010F7",
INIT_21 => X"5D556AA00FFAE95555AAFFE8A00552EBFE00F7D17FF45F7FFFFF55AA80155FF0",
INIT_22 => X"AAAAAA8B55F7D140010552E821EFAAAABDF555555555EFAAFFFDFEFAAAAAAB45",
INIT_23 => X"45557BE8A00AAAE955450055421FFFFFBC0010AAD5574BA557FFDFFF5504000A",
INIT_24 => X"FFFF7FBEAA00002EAAAAA082EA8A00002AA8A10F78402155AA8028A00A2D57FF",
INIT_25 => X"75D7000000000000000000000000000000000000000000000557BFDFFF55003D",
INIT_26 => X"FAE105D556AA10410E17555080E000280071E8A00EB8E3FE10F7AEBAFFF080A1",
INIT_27 => X"EA8AAA5571C2000FF8A17400557FC015514555757DFF8E175C7A2AAAAA82A2F1",
INIT_28 => X"FFF8F7DB68A105D71C7BFFF55FFA095482B6A49256DEB84104BAFFD1525FF492",
INIT_29 => X"AF1FFFD7AAAAAFB7D495F6AA10E3AE90555A2FBE8A38492ABDE10EBDF7AF6DE3",
INIT_2A => X"5571FDFEF550E00082B6A0AFB55F7D1420104124821D7AAA0BDF6D415B575D7A",
INIT_2B => X"DA2842FA00B6D578F6D557FFDA00A2AE9756D145B401FFFFFFC7010BEDF524AA",
INIT_2C => X"00497BFAFFF49003AFEFEBFBEAA001C2EA8A821C2EAAA001C2EA8A00F7800017",
INIT_2D => X"E00F7AEAABEF082E955450000000000000000000000000000000000000000000",
INIT_2E => X"7555A2AEA8A10AAD568A00555168A10002E9754D082E820BA08556AA00AAAABF",
INIT_2F => X"000AAFFD1401E7082EAAABA5D5140010F7AE974105D7BC21555D51575EFFFAA9",
INIT_30 => X"ABFE00AAFBEABFFAAFBEABFFF7AA80145557BFDF55F78017400F780001FFAA84",
INIT_31 => X"843FFFF007BD5555AAD57DF55AAAEBDFEF007BE8A10AAAE8215DA2FFE8ABA082",
INIT_32 => X"7FBD7400F7FBC00BA55557DFF75D2E82010F7843DF45FFD540000000402145AA",
INIT_33 => X"5D2AAAA10F780021FFA2803DE10FFD16ABFF5D7BFDE10AAAA975FF5D7BC21EFF",
INIT_34 => X"0000000000000000000007FE8BFF080028BFFAAFFEAA105D2EAAA005D2AAAA18",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000400000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000006",
INIT_01 => X"000009801830084C182060000C104268413C0A61590001D90213C10008110200",
INIT_02 => X"680108200010000054400C000080000041000000010002400800800009082011",
INIT_03 => X"0008000004002040000200100000000042800504488000103081880008C00000",
INIT_04 => X"00005042802A82100010030018000010000040C0100040140080040800003100",
INIT_05 => X"2000200400245001012100006002082000000000004000002010000040002000",
INIT_06 => X"2320400004040040144A7D000180020101000009808000000800001008210000",
INIT_07 => X"6100000021808000940800001800010200018B20206C01020200002441223C12",
INIT_08 => X"184010110120000004000000000061F000000244000081180004400000400000",
INIT_09 => X"4111002100040010008528820005100000900280000001000550860020002800",
INIT_0A => X"0080200520B23204000116404470900100402000000100242048025481024010",
INIT_0B => X"400000115040008002200000048034000002000000010712000000800F08A505",
INIT_0C => X"0000410004000041000400004100020000208201000000200404840284500016",
INIT_0D => X"00000120040000080000900201A0021924600088000000100100041000410004",
INIT_0E => X"60002000120002121C99024A00A14650A328519428651900142000000200A008",
INIT_0F => X"0000A20010200900000001400008200900000001400000001424008208041001",
INIT_10 => X"000002400820090000000140000820090000000140000A800000000000000000",
INIT_11 => X"0000000000000001500012000200800000000000000C10008400080200000000",
INIT_12 => X"0000000480004800002040000001000400000000000000004800010002800000",
INIT_13 => X"8041000000002401F80000000000000000025000274020800000001205D00808",
INIT_14 => X"004020000000000002900009AB00200800000000000012BA010100000000902E",
INIT_15 => X"652035000104000000000000001040100009BA000000000000000005400023B8",
INIT_16 => X"19028CA8D06540144C26832A1B0004000020024048400000090032A000000010",
INIT_17 => X"9425094250942509425094250942509425094250942509425094251946519465",
INIT_18 => X"4250942509425094250942519465194651946519465194651946519465194651",
INIT_19 => X"0800000000000000001465194651946519465194651946519425094250942509",
INIT_1A => X"34D34D1285B080201C92410480AB9A26667A46F345448020082E1C712A054008",
INIT_1B => X"1A0D068341A0D06834514514514514514514514514514514514514514D34D34D",
INIT_1C => X"2B60D069349A0D068341A4D268341A4D268341A0D069349A0D069349A0D06834",
INIT_1D => X"0000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF829",
INIT_1E => X"0155FFAAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA0000000000000",
INIT_1F => X"FBFDFFFA2AEBDE00AAFBEAABA080000000087BEAA10F7803DE00FFAEBFFFF080",
INIT_20 => X"780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555087BFDE00A2FBD7400F7",
INIT_21 => X"5D7FC2145005155555557BE8BEF007FFDEAAAAD1555EF0055401FFF7AEAAA10F",
INIT_22 => X"A5D2AA8A10F7AA974AA082E80010A2AAAAA10552AA8AAA557FC0010F78015410",
INIT_23 => X"45002EAAABA087BFDF45F7AA974AAAAAA97555F784174BAF7D5555FFF780154A",
INIT_24 => X"E00F7D17FF45F7FFFFF55AA80155FF080400145FFFBEAABAF7D17FEBAA2AEBDF",
INIT_25 => X"8A92000000000000000000000000000000000000000000000AAFFE8A00552EBF",
INIT_26 => X"3FE10F7AEBAFFF080A175D7BEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E",
INIT_27 => X"1FFE00A2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92080E000280071E8A00EB8E",
INIT_28 => X"5B451D7FFAAA8A38FF8E175C7A2AAAAA82A2F1FAE105D556AA10410E17555087",
INIT_29 => X"571C2000FF8A17400557FC015514555757D5D71E8BEF147BFAE82A2DB555C71C",
INIT_2A => X"FFD1525FFFF84174BA5D20AAA00E3AA904BA142A87010A2AEADA38492EA8AAA5",
INIT_2B => X"2FFD57DEBAAAA0BFF7D0024ADA921C7BFFF55FFA095482B6A49256DEB84104BA",
INIT_2C => X"00A2FBE8A38492ABDE10EBDF7AF6DE3FFF8F7DB68A105D7000400155FFFBEDA8",
INIT_2D => X"B55FFAABDFEFF7D16AA000000000000000000000000000000000000000000000",
INIT_2E => X"20BA08556AA00AAAABFE00F7AEAABEF082E95545F7D568BEF080402000F7AAA8",
INIT_2F => X"68A10002E9754D00517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00082E8",
INIT_30 => X"FE8A10AAFFD55555D7FD5555FFAAA8AAAFFAA97555A2AEA8A10AAD568A005551",
INIT_31 => X"AEBDEAA082EAAABA5D5140010F7AE974105D7BC21555D51575EF555568BEF5D7",
INIT_32 => X"780001FFAA84000AAFFD1401E7FF80174AA5D0028A00AAAE800AA552A97400A2",
INIT_33 => X"080002145F7FBFFE00FFD17FEAAA2803DFEF08043FE00557BFDF55F78017400F",
INIT_34 => X"0000000000000000000A2FFE8ABA082ABFE00AAFBEABFFAAFBEABFFF7AA80145",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000800000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A14009821830284D182060000C10426840000000080000080200080000510204",
INIT_02 => X"0801080200100000046558040080000041000000002402400800000009008010",
INIT_03 => X"00020201040000D0842242024210810802006400088000003080054288C10000",
INIT_04 => X"0000400088020000003020002000001002A0E881108032100002000800203040",
INIT_05 => X"200000040000004924040108022000201000012800400010001081C040402000",
INIT_06 => X"030040040404804100006D2002A002012120004CC08125410200082308290000",
INIT_07 => X"2181020421408000940820001800010200018920206C01020200002440003C00",
INIT_08 => X"084010110120018004000000000021F020408264000000080004400800400000",
INIT_09 => X"511110010100008210010802004404230A000888400809000010042002002800",
INIT_0A => X"0000200000C04204000116404460910100082000040100240000000000004010",
INIT_0B => X"0AE22291404020902005002010000420A0200000400414684920410420200000",
INIT_0C => X"1120001200012001120011200011000090008840221000240484110000F05044",
INIT_0D => X"000803004C150100088480000980020000050001011890008011000120011200",
INIT_0E => X"000060001000020010010248040200010000800241000008009042404003E0BC",
INIT_0F => X"0080A00010202800000001402008202800000001402000000026008208041001",
INIT_10 => X"0000034008202100000001402008202100000001402002800000800000000000",
INIT_11 => X"8000000000000081400012000300000000000000008C10008400081000000000",
INIT_12 => X"8000000680001040002040000001000100000000000000004810000002800000",
INIT_13 => X"0001200000003408000004000000000040027000200020100000001A00000800",
INIT_14 => X"004010000000000042B00001000020800000000000801200000110000000D000",
INIT_15 => X"0000000001000100000000000010C030000100000200000000000105C0002000",
INIT_16 => X"03700080022100404D26A42EA01004002022000080000000018032A000A00010",
INIT_17 => X"0040100401004010040100401004010040100401004010040100400000000200",
INIT_18 => X"0000000000000000000000010040100401004010040100401004010040100401",
INIT_19 => X"0800000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"8A28A28D532A0CCC2A28A28A7AA344854A07F069CB8930AFD6A1AAA902A14148",
INIT_1B => X"6532994CA6532994CA28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A2",
INIT_1C => X"CC772B94CA6532994CA6572B95CAE532994CA6532995CAE572B94CA6532994CA",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF831",
INIT_1E => X"FEAABA007FC2155F7D155545AA80001EFAAFBEAB45557FFDE100000000000000",
INIT_1F => X"8000010FFFBE8BFFF78402155AAFBE8B45002A974AAAA803DFFFAA843DF45FFF",
INIT_20 => X"80000000087BEAA10F7803DE00FFAEBFFFF0800155FF00042AB55FFD168B55AA",
INIT_21 => X"A2AEBDE00AAFBEAABAA2FFD741055003DFEFF7AA801FFAAD16AABA002ABDE100",
INIT_22 => X"05555555EFF7FBC0145F78028A00A2D142155087BFDE00A2FBD7400F7FBFDFFF",
INIT_23 => X"FFF7AEBDEBAF780155EFAAAEA8ABAAAFBFDE0055556AA005D0415555007FD741",
INIT_24 => X"EAAAAD1555EF0055401FFF7AEAAA105D042ABFF5D556AB55AAD168ABA002A975",
INIT_25 => X"8E00000000000000000000000000000000000000000000000557BE8BEF007FFD",
INIT_26 => X"38FC7BE8A3DF7DF7F5E8A92007BC217DEBDB55555AA8E071D7AAFBEFB455D71F",
INIT_27 => X"42AB7DEBDB6DB55BE8E05000EBFFE8BC7E38E07145BEF1E8B6D002090482B68E",
INIT_28 => X"D16FA82142EB8E00080E000280071E8A00EB8E3FE10F7AEBAFFF080A175D7000",
INIT_29 => X"2FBD0400FFF5FDFC7B6A0BDE38B6F5E8A92B6FBD5410490A3DFD7F7A4821D7A2",
INIT_2A => X"410E175550071D54104951555D7EBF5C5155E3842AA00BED1421450871FFE00A",
INIT_2B => X"5BED16FA820820955EFE3AEBDEAAFF8E175C7A2AAAAA82A2F1FAE105D556AA10",
INIT_2C => X"005D71E8BEF147BFAE82A2DB555C71C5B451D7FFAAA8A38410E2ABD749516FB5",
INIT_2D => X"555A2FBFDF455D556AA000000000000000000000000000000000000000000000",
INIT_2E => X"8BEF080402000F7AAA8B55FFAABDFEFF7D16AA00087FC01EFA2FFD7545AAAE97",
INIT_2F => X"AABEF082E9554500042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D56",
INIT_30 => X"EBFF45F78400155A2D57FE00552EA8A00082E820BA08556AA00AAAABFE00F7AE",
INIT_31 => X"D54214500517DE00A2FFC2000F7D17FF55FF803FEAAFFD16AA00FFFBD5400082",
INIT_32 => X"AD568A00555168A10002E9754D085155410085557555AAD557555A2802AA10FF",
INIT_33 => X"002AAAB4508557DF55F7D17FE000804155FFAAAABDEAAFFAA97555A2AEA8A10A",
INIT_34 => X"0000000000000000000555568BEF5D7FE8A10AAFFD55555D7FD5555FFAAA8AAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000008FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400986B830284D1820E0000C3642484000000008000008820009080A512220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"00080D4912E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"000048048002400048150300100002504230C8D9109032100020160880223000",
INIT_05 => X"220004440040080142020015001004A01200012840440000B01088C0005C2400",
INIT_06 => X"431018040014804920906C74B320020121210045408165445220082008211002",
INIT_07 => X"A5B1220421408004A56E840008B90D0200018B60A0650D450FC800644A0438A0",
INIT_08 => X"485816170760268E04000000000323F42C50826490640D28088445B0E0419003",
INIT_09 => X"41F1654100000818128728820024002B3B01AC9540080824CA13008820A02800",
INIT_0A => X"0000203600E06204000116C14474A3650048CE64E40100260048025481024810",
INIT_0B => X"08C32E915D9C208070042420180D24C8802000284007126A4D21262C20200404",
INIT_0C => X"31CA821CA831CA831CA821CA83165410E541085102000024040490A000D01056",
INIT_0D => X"812203360410110A4000840E3180021040465501011934A005101431CA821CA8",
INIT_0E => X"60006000101004A01811064B050204810240812241280D00200A08044290A088",
INIT_0F => X"482A01AAEC3602330CD2A02952DC3502330CB4A0318B41400024008208041011",
INIT_10 => X"0144C0155C3502330CD2A02952DC3602330CB4A0318B5600C587149B6D0141B0",
INIT_11 => X"083B6A51005956308D1E8202C436375908AA840AD4513437640F15245B455163",
INIT_12 => X"62F47B2872400044959BC42B1060F0D036B80B548523136C158878D8FE04E587",
INIT_13 => X"0A2699AAA3794392000D81852B0A050C224180062085134CD1719564E020C670",
INIT_14 => X"C50500D94C8121713C02B555101C90705D71009604140C0418CE0C378F0B2701",
INIT_15 => X"828E024D8C50965A40821568A06113801505010334AA73AA0666DAC20AD57400",
INIT_16 => X"123408C0822040544D248604B2100400100084008001D0113920060CDC06A27C",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"0080200802008020080200812048120481204812048120481204812048120481",
INIT_19 => X"0000000000000000002008020080200802008020080200802008020080200802",
INIT_1A => X"2082082815220A4A380000002A8313044020C0605885026853A1082100A00142",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000008208208",
INIT_1C => X"F070000000000000100800000000000000000004020000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF801",
INIT_1E => X"FFDE10082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA0000000000000",
INIT_1F => X"2A801FFF7FFE8A10A28000000007FC2155F7D155545AA80001EFAAFBEAB45557",
INIT_20 => X"AFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABAA2AEBFF45FFAEBFEAA00",
INIT_21 => X"FFFBE8BFFF78402155AAD155555A28428BFF002ABDE00A2AABFE10082ABFFEFA",
INIT_22 => X"5557FC2010002A80010A2842AAAA007BFFF4500042AB55FFD168B55AA8000010",
INIT_23 => X"EFFFD540000080000000087BEAA10F7803DE00FFAEBFFFF0800155FF00557FF4",
INIT_24 => X"FEFF7AA801FFAAD16AABA002ABDE10A2D168A10A284021FF5D00154BAF7FBE8B",
INIT_25 => X"70AA000000000000000000000000000000000000000000000A2FFD741055003D",
INIT_26 => X"071D7AAFBEFB455D71F8E00002EBDF6D005B78F7D142ABDFC7F78E3FE28B6840",
INIT_27 => X"EBFF7DEBA0BDEAA1C2A801C7E3FFEFA10B68407038007BC217DEBDB55555AA8E",
INIT_28 => X"AAB8E280820B8FEFBEF1E8B6D002090482B68E38FC7BE8A3DF7DF7F5E8A92BEA",
INIT_29 => X"BDB6DB55BE8E05000EBFFE8BC7E38E07145B6D15756DA28A28BFF082ABAE10B6",
INIT_2A => X"080A175D708517DF7D497BC5028142A87000A28A2AA92007FF8F7D00042AB7DE",
INIT_2B => X"F5D0A10482FFFFEFBC7E3DF42028080E000280071E8A00EB8E3FE10F7AEBAFFF",
INIT_2C => X"00B6FBD5410490A3DFD7F7A4821D7A2D16FA82142EB8E00B6DB6AA28A280001F",
INIT_2D => X"F55F7AABDEAAF784154BA0000000000000000000000000000000000000000000",
INIT_2E => X"01EFA2FFD7545AAAE97555A2FBFDF455D556AA00082EBFFEF007BE8BFF5D2ABD",
INIT_2F => X"BDFEFF7D16AA00FFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BA087FC",
INIT_30 => X"AA8BFF002AAAA00FFAAA8AAA080028BFFF7D568BEF080402000F7AAA8B55FFAA",
INIT_31 => X"7FEABFF00042ABFFA2FFFFF45F7AE97400AAFFE8B45AAAA95545F7D5555FFAAA",
INIT_32 => X"AAABFE00F7AEAABEF082E9554508557DFFF007BD54BA5D2E95400A2AEA8A0000",
INIT_33 => X"FFFFE8AAAAA80001FF5D2E82000F7FFFFF45AAFFC20BA082E820BA08556AA00A",
INIT_34 => X"0000000000000000000FFFBD5400082EBFF45F78400155A2D57FE00552EA8A00",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000800000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702484000000008000008820009280A553231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"421A0A0012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"02004000890200001837830011998C31C09060DC104000102002140900003548",
INIT_05 => X"240000C400000001E404001F064000A00800000020480010A4100100001C2000",
INIT_06 => X"0300D800C1960C4400006E10B900020181840001008040057840001308212000",
INIT_07 => X"652428112180C03E8E5A2C800A3F018200418927E06686450FF8006460003A00",
INIT_08 => X"9840903525281D4F460409000000E3F08D1202C5C26A0719CC96CC7BF4629900",
INIT_09 => X"491175E10000041000C52882008600843001E09F0000002CF810200022302800",
INIT_0A => X"00002000030003040081164FC469227D2008CFE09A8180248009021091004810",
INIT_0B => X"00010C13499F01B33A00ACC0000F04F800000011800000000000433800000000",
INIT_0C => X"20CBC20CBC30CBC20CBC20CBC3065E1865E1000100000820040482B280504016",
INIT_0D => X"E7F3F01F40401C17E800C7FF3B80020000035780460124F16F06BC20CBC30CBC",
INIT_0E => X"00002200004005002001408400000000000000000000053A4096F80705FA0201",
INIT_0F => X"7B2C53F2FC16691DB587201EDDF4162B1DB527201EDDC46070241001000200F5",
INIT_10 => X"01D5CC9794162B1DB587201EDDF416691DB527201EDDD884272592D6246FC1B1",
INIT_11 => X"8E995D5A825DBA569F9FF02547068618CD3CC45B7863AE7EC00D4B122A67DF2A",
INIT_12 => X"CA5C33717461C045B5B182019473D19D7CCD856106F31A683621BDFC28800725",
INIT_13 => X"0A652CC8E3538BBA01624E51AA6C0469AC5493F5688532966471A9C5F6208C6C",
INIT_14 => X"41E1F5759001B4AA1853E6D5144AA9C914C8608D2724A4C4118D992B866E2FB1",
INIT_15 => X"825682D4A36C0B0B4B85112B2C4A05D3E6D5051893335EB0072AA85A4F9B7400",
INIT_16 => X"00800000082100544D248020000004001DC0800000010E7F70171401DE07EAD9",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0401004010040100401004000000000000000000000000000000000000000000",
INIT_19 => X"0800000000000000000040100401004010040100401004010040100401004010",
INIT_1A => X"249249120780800016A28A288028DCA30444409B054A88C5890486582A210108",
INIT_1B => X"32190C86432190C8641041041041041041041041041041041041041049249249",
INIT_1C => X"007592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2592C864",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF83E",
INIT_1E => X"0000AAAA843FE0008557DFFF0800020105D557FEAA00557DE100000000000000",
INIT_1F => X"AA8200000557DFFFF7AA80000082ABDF5508557DF45002ABDFFFF7803DE10AA8",
INIT_20 => X"07FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AAD5420000051555FFA2",
INIT_21 => X"F7FFE8A10A28000000A2D155410F7FFFFEBA08003FE00082AA8AAAAAFFC00BA0",
INIT_22 => X"05D2ABFE10A2AABFE1055516ABEF5D517DEAAA2AEBFF45FFAEBFEAA002A801FF",
INIT_23 => X"FFF7AA82155AAFBE8B45002A974AAAA803DFFFAA843DF45FFFFEAABA000028A1",
INIT_24 => X"BFF002ABDE00A2AABFE10082ABFFEF085542000000417555002A820AA08557DF",
INIT_25 => X"DE10000000000000000000000000000000000000000000000AAD155555A28428",
INIT_26 => X"BDFC7F78E3FE28B684070AABE803AE38145B78FD7000005010495B7AE921C517",
INIT_27 => X"547038145B505FFB6A487000005F7AFD7F7A482038002EBDF6D005B78F7D142A",
INIT_28 => X"2EAAAAAB6F5C2082007BC217DEBDB55555AA8E071D7AAFBEFB455D71F8E00BED",
INIT_29 => X"BA0BDEAA1C2A801C7E3FFEFA10B68407038B6D550428FFF1FDE821C003FE001C",
INIT_2A => X"F7F5E8A9200002FA285D20BDE28A2A4B8E10555B68BEF5D517DEAABEAEBFF7DE",
INIT_2B => X"5142082082005F7DFD7F7A482155BEF1E8B6D002090482B68E38FC7BE8A3DF7D",
INIT_2C => X"00B6D15756DA28A28BFF082ABAE10B6AAB8E280820B8FEF085F4703814001055",
INIT_2D => X"410007FEAA0055517DE000000000000000000000000000000000000000000000",
INIT_2E => X"FFEF007BE8BFF5D2ABDF55F7AABDEAAF784154BAF7802AABA5D7FEAB45080015",
INIT_2F => X"FDF455D556AA00F7D1554BA5D7BC01FFFF8015410007FEAB45F780020BA082EB",
INIT_30 => X"57FE005D043FE10552EAAAAAFFD140000087FC01EFA2FFD7545AAAE97555A2FB",
INIT_31 => X"557DEBAFFAEBFFEFAA803DEBA5D2E82155A2FBFDE00FF84154BAF7D1400BAFFD",
INIT_32 => X"7AAA8B55FFAABDFEFF7D16AA0008003FEBA55003DEBAA28428A105D7FEABEF55",
INIT_33 => X"087BD54AA550402145550000010087FFFF45F78402145F7D568BEF080402000F",
INIT_34 => X"0000000000000000000F7D5555FFAAAAA8BFF002AAAA00FFAAA8AAA080028BFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042604001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00020201926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"00104884880A4400403000004800027102A0E88110D83210642EA809C0203040",
INIT_05 => X"27000004004828032646000826080C201A008128044E00754010C9C192D82400",
INIT_06 => X"43000004080480492A946CE10320020121258044408125410270082308213800",
INIT_07 => X"A581424525408000AE2AA8002BC00D020003896020658FC4030000246E543AE5",
INIT_08 => X"4840101107200B80040210000002ABF02450A264002C80080004416800419000",
INIT_09 => X"4B531001000008001041080200B660E30B200C8840080A920651020002802800",
INIT_0A => X"0000203240E46204000516C04468C10100540034AC0100259001004010025010",
INIT_0B => X"04462E91440020905200A42209002420002800284002026A4D21758400000000",
INIT_0C => X"10000000000000010000000000000008000000000000002004040AA080504004",
INIT_0D => X"00000360401021280800E4000B800610C8410000A11210000000001000000000",
INIT_0E => X"6000600040D045E4195104D5854284A14250A12A512A8808289840084A020080",
INIT_0F => X"9E07A80948354B6E68982167061037496E683821670620681024000000000008",
INIT_10 => X"10B456587037496E689821670610354B6E6838216706220431961CA985D48094",
INIT_11 => X"186A91674011CE61403562274AA49CD594CF00039C7C414B6509DA22652138E5",
INIT_12 => X"3014780CC8604040424A5323845932E620295879818170304B2F5002C2043196",
INIT_13 => X"654B9104A328665603148895D44E0251142B42A3D8B2A5C8825194328A2E6A98",
INIT_14 => X"A6C6A465AA0091482382B17614F2202858EE300991415B45CD5306028F019451",
INIT_15 => X"08DC8047F17D1C7C3C02128E587D6A02B17605A130A4E8BF002258850AC5DC06",
INIT_16 => X"123508508220808048260604B2100C00022084809000D000393722A14000052E",
INIT_17 => X"284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A",
INIT_18 => X"84A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1",
INIT_19 => X"000000000000000000284A1284A1284A1284A1284A1284A1284A1284A1284A12",
INIT_1A => X"BAEBAEBFF6FEFEFEEEAAAAAAFBF7DDF77F9FBEFBFF9F3F0FDFCFBEFBF1228154",
INIT_1B => X"FD7EBF5FAFD7EBF5FAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAE",
INIT_1C => X"0077EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FA",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"57DE10AAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF0000000000000",
INIT_1F => X"7BEAB45552E80155AA802AB45AA843FE0008557DFFF0800020105D557FEAA005",
INIT_20 => X"82ABDF5508557DF45002ABDFFFF7803DE10AA80000AA087BD75EF087FFFFEF55",
INIT_21 => X"00557DFFFF7AA80000AAD1420AA087BD7555FFD168AAAFFAE820AA5D55575550",
INIT_22 => X"FA2FBD7545FFD157555085140010F7AEAABFFAAD5420000051555FFA2AA82000",
INIT_23 => X"BAFFAAAAB45007FC2155F7D155545AA80001EFAAFBEAB45557FFDE10AAAEA8BF",
INIT_24 => X"EBA08003FE00082AA8AAAAAFFC00BA00002AAAAF7D5574BA557BE8A10A284154",
INIT_25 => X"ABD7000000000000000000000000000000000000000000000A2D155410F7FFFF",
INIT_26 => X"05010495B7AE921C517DE10A2DB50482147FFAF554971D0492E3F1C71C7BE8A2",
INIT_27 => X"1D25D7007FFAFD7497BE8B5555208217DBE8A2AB45BE803AE38145B78FD70000",
INIT_28 => X"A4870BA555F5056D002EBDF6D005B78F7D142ABDFC7F78E3FE28B684070AA1C7",
INIT_29 => X"45B505FFB6A487000005F7AFD7F7A482038AADF47092147FD257DFFD568A82FF",
INIT_2A => X"5D71F8E00A2A0ADBC7A2FFD257DE3DF52555085142000FFAAAFBFFBED5470381",
INIT_2B => X"24171EAA10B680124BAFFAAAFB45007BC217DEBDB55555AA8E071D7AAFBEFB45",
INIT_2C => X"00B6D550428FFF1FDE821C003FE001C2EAAAAAB6F5C20821C002AA92FFDF5748",
INIT_2D => X"010AAD157545F7AEA8B550000000000000000000000000000000000000000000",
INIT_2E => X"AABA5D7FEAB45080015410007FEAA0055517DE00A2FFC00105D7BE8B55085142",
INIT_2F => X"BDEAAF784154BA5D5140145007BE8B55087BEAB555D04001EFF7AAA8B55F7802",
INIT_30 => X"FC21EFFFD16AA10FF80174AA557FC21EF082EBFFEF007BE8BFF5D2ABDF55F7AA",
INIT_31 => X"AEBFFEFF7D1554BA5D7BC01FFFF8015410007FEAB45F780020BAA2FFD54105D7",
INIT_32 => X"AAE97555A2FBFDF455D556AA00A2803FF45AAFFC21EFAAFBC0155085540000FF",
INIT_33 => X"5D042AA00F7FBD5410085568A10FF80020AAFFAABFF55087FC01EFA2FFD7545A",
INIT_34 => X"0000000000000000000F7D1400BAFFD57FE005D043FE10552EAAAAAFFD140000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000CFFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"0002074F200904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000480488024000403000000000001002A0E881108032100002000800203040",
INIT_05 => X"200000040040080126060008020000201000012800400010001081C000402000",
INIT_06 => X"430000040004804920906C200220020121200044408125410200082308210000",
INIT_07 => X"A5A14285A15080008768A80008000D0200018B202067AF100A00002442043820",
INIT_08 => X"4850101105205380040000000000A7F42840A264920406080004400A00409002",
INIT_09 => X"411110010000080010010802000400230B000C88400808000211000002002800",
INIT_0A => X"0000203200E0620400011640446DA101004000002C0100240000000000004010",
INIT_0B => X"00422291400020900000002008002420002000004000026A4920410400000000",
INIT_0C => X"0000000000100000000000000100000000000000000000200404000000504004",
INIT_0D => X"0000022040100108080080000B80021040410000011010000000001000010000",
INIT_0E => X"0000600000000020181100400502048102408122412808082098400042020080",
INIT_0F => X"0040A100A42008000161C140000420080001C1C1400003201024000000000000",
INIT_10 => X"00022260042001000161C140000420010001C1C140001604E8084341CBA34048",
INIT_11 => X"2580E2B8802201014800C220A21829A302F1C024010C001124020C8C1A8A0396",
INIT_12 => X"0CA000048228404401004418012787124648157780120B8678C000801E04E808",
INIT_13 => X"072D04730000241000CB1325E78E0186030240000083B602398000120024ACA6",
INIT_14 => X"EF6F4163C480481506800004000CFD55196CB012481812049495C19400009001",
INIT_15 => X"800108B8FB61A0401200845594965000000400568D0CFB780055060500001001",
INIT_16 => X"123408408220000048240604B210040000008400800B0000090022A140068248",
INIT_17 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_18 => X"0481204812048120481204812048120481204812048120481204812048120481",
INIT_19 => X"0000000000000000002048120481204812048120481204812048120481204812",
INIT_1A => X"9E79E79FF3BEEEEEFE79E79EFAABCDA72E47F87BDF4EBAE7CFAFBEFB28200140",
INIT_1B => X"7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"FF83F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF83F",
INIT_1E => X"02ABEFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA0000000000000",
INIT_1F => X"AE955455500155EF0804155EFAAD5554BA087FFFF55557BD54AAF7FBC01FFA28",
INIT_20 => X"A843FE0008557DFFF0800020105D557FEAA00557DE10A2AA801FFA28402000AA",
INIT_21 => X"552E80155AA802AB4500516AA00A2AE800BAFFFFC20BAF7AEA8B45080417400A",
INIT_22 => X"AA28402010A2843FEBAFFFBD7410A2D168BFF087BD75EF087FFFFEF557BEAB45",
INIT_23 => X"EF00043FEAA082ABDF5508557DF45002ABDFFFF7803DE10AA80000AA005568AB",
INIT_24 => X"555FFD168AAAFFAE820AA5D5557555002E80155A280000005D7FFDF4555517DF",
INIT_25 => X"0092000000000000000000000000000000000000000000000AAD1420AA087BD7",
INIT_26 => X"D0492E3F1C71C7BE8A2ABD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB4",
INIT_27 => X"E851FFB68402038AAAA955554900105FF0800175D7A2DB50482147FFAF554971",
INIT_28 => X"AAADB6D080A12410BE803AE38145B78FD7000005010495B7AE921C517DE10A2A",
INIT_29 => X"07FFAFD7497BE8B5555208217DBE8A2AB451C556FA00A2A0800BAE3F1C0092EB",
INIT_2A => X"B684070AA00516DABAA28402038B6803DE82F7F5D5410A2D568BC71C71D25D70",
INIT_2B => X"05D7FF8F455D5F78FD7000E3FEAA002EBDF6D005B78F7D142ABDFC7F78E3FE28",
INIT_2C => X"00AADF47092147FD257DFFD568A82FFA4870BA555F5056D002A80155B6800001",
INIT_2D => X"145002AA8AAAAAFFC20000000000000000000000000000000000000000000000",
INIT_2E => X"00105D7BE8B55085142010AAD157545F7AEA8B55A2FBFFF55FF84000AAAAFBC0",
INIT_2F => X"EAA0055517DE00A2AA955FFFF80020BAAAAA975450800001EF080417555A2FFC",
INIT_30 => X"0020BAAAD140000A2AEBFFEF082A82010F7802AABA5D7FEAB45080015410007F",
INIT_31 => X"D56AB455D5140145007BE8B55087BEAB555D04001EFF7AAA8B555D557FE00A28",
INIT_32 => X"D2ABDF55F7AABDEAAF784154BA08557FEAAA284000AAFF803DE00FFD557400AA",
INIT_33 => X"082A80145F780020105D7BEAB45557BE8B45082EBFEBA082EBFFEF007BE8BFF5",
INIT_34 => X"0000000000000000000A2FFD54105D7FC21EFFFD16AA10FF80174AA557FC21EF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000100000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"000440009282000001100000000000100220C8811080321000000228002A3000",
INIT_05 => X"200014C40000000100000000005C04A01000012A64400000145080C000422000",
INIT_06 => X"031042040804804100006EE4032002012120005540812540020008600831000A",
INIT_07 => X"21912244A14080008408880008000D0200018920206563000200002440003800",
INIT_08 => X"48501415032000800406180000002DF024408264000000080004400000430800",
INIT_09 => X"411100110000000010010802000400230A000880400808000450200000B02800",
INIT_0A => X"0000203000C042040001164044608101000000007C0100240000000000005810",
INIT_0B => X"0042229140002080000000200000040000200000400000684920000400000000",
INIT_0C => X"1000010000000000000000000100000800008000000000200404000010500004",
INIT_0D => X"00000260001001280000C4000300020000000000011010000000001000010000",
INIT_0E => X"400060000000000010010040040000000000000201000000000000004A000080",
INIT_0F => X"0000000000202100000000000000202100000000000004600024000000000008",
INIT_10 => X"0000000000202800000000000000202800000000000002000000800000000000",
INIT_11 => X"8000000000000000000002000100800000000000000000000400001200000000",
INIT_12 => X"80000000006000400080C0000000000D08120280000000000000000002000000",
INIT_13 => X"0040200000000010000004020010000000000000008000900000000000200008",
INIT_14 => X"0000308801400000000000040000008822110000000000040100100000000001",
INIT_15 => X"0000000004840717050000000000000000040000020000000000000000001000",
INIT_16 => X"023000000220000048240404A010040000008000000000000000020C40000008",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000200140",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"1420BAFF8000010082A954BA00003DFEF085155400F78428BEF0000000000000",
INIT_1F => X"843DE00AA8015400FF84001EFA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD",
INIT_20 => X"AD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEFF7AE95555A2FBE8BEFA2",
INIT_21 => X"5500155EF0804155EFFFFBE8BFF0800174AA557BFDE10A2FBEAB45F7D56AABAA",
INIT_22 => X"AA2D16AB55FFD568BEF087FE8A1055003FE00A2AA801FFA28402000AAAE95545",
INIT_23 => X"BA5D0015545AA843FE0008557DFFF0800020105D557FEAA00557DE10F7D1574A",
INIT_24 => X"0BAFFFFC20BAF7AEA8B45080417400FFFFC2145080015400AA802AA00AAAE800",
INIT_25 => X"DBFF00000000000000000000000000000000000000000000000516AA00A2AE80",
INIT_26 => X"50555412AA8ABAAADB40092E38E070280024904AA1C0438FD7005150438F78A2",
INIT_27 => X"A9257DA2FFE8BC7BE8E38E10A28017400E38A051FFA2FFEDB55B6A080038E3DB",
INIT_28 => X"FBEDB6DF7D16AABAA2DB50482147FFAF554971D0492E3F1C71C7BE8A2ABD7E3A",
INIT_29 => X"68402038AAAA955554900105FF0800175D7E3FFEFBD70000124AA557FFDE10A2",
INIT_2A => X"1C517DE10FFDF50482A2DB6AB45FFD56DBD7087BEAA38410038E38A2AE851FFB",
INIT_2B => X"0BE8E28A10AAA085082550A1057DBE803AE38145B78FD7000005010495B7AE92",
INIT_2C => X"001C556FA00A2A0800BAE3F1C0092EBAAADB6D080A12410FFF1C017D14041040",
INIT_2D => X"B550855400AAF7AEBDFEF0000000000000000000000000000000000000000000",
INIT_2E => X"FF55FF84000AAAAFBC0145002AA8AAAAAFFC2000AAAA974AA0800020BA550028",
INIT_2F => X"57545F7AEA8B55AAAE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EFA2FBF",
INIT_30 => X"4020AA557BFFE10A2FFFFFEFF7D568ABAA2FFC00105D7BE8B55085142010AAD1",
INIT_31 => X"002AAAAA2AA955FFFF80020BAAAAA975450800001EF080417555AAFFFDF45080",
INIT_32 => X"80015410007FEAA0055517DE00FFFBC2000AAFBE8B55F7D17DF45007FE8AAA08",
INIT_33 => X"FFD5421EF5D0000010F7AAA8A10AA8017400552A801EFF7802AABA5D7FEAB450",
INIT_34 => X"00000000000000000005D557FE00A280020BAAAD140000A2AEBFFEF082A82010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000C00000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"0202115002BB10080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"2FE962000017102918900948514522CE09200C0D590569398ADBF8CC1E50E480",
INIT_05 => X"F05EA11E5600006B0800000038814B72A15B71D412E0AFD9C2990DA56FF0B55A",
INIT_06 => X"0640044150C025A0000000901A054F2C0A8030140BCC0460050690A95C8383D0",
INIT_07 => X"288500102F85203E8010D0AA9BC4800015001219D0550077373CAA8040006800",
INIT_08 => X"2064193920A2004B51400001414091EAA14881C0002701881B120203B7A80120",
INIT_09 => X"0409A02D965965200100104F2B00822512000000231520A024400800000ACCAA",
INIT_0A => X"0004B240028000342A00002FE00A3A1F06E649C005514AC40C082050010222D9",
INIT_0B => X"000A448C0082024AE50064B44000000000002A296AA000604838001980000000",
INIT_0C => X"044000440004400044000440004200022000200014808A02004200E540480212",
INIT_0D => X"0A80A5C8000102ED00440630004AD32400004000D58460018F6D3D8440004400",
INIT_0E => X"12AA28AA890BA00000024800480000000000000200802151025062C0BB400014",
INIT_0F => X"54E11C596A64003195933741477264003195555B418687E35836020814004049",
INIT_10 => X"99CF47DCB264003195933741597264003195555B4198843940076D296D0031F5",
INIT_11 => X"58486A556489347FE5F409CBC1362510695B6288743123C95251852041CD50A4",
INIT_12 => X"EAE2992046EB70026486035600CEC45CBCA809654B48163CCC895E1E043D4007",
INIT_13 => X"3A242DEA151848302BFD6D522B10C7EC71F6C1DB071D1216E078C4C1B1C74424",
INIT_14 => X"DAAABC982BE22267A2E2E4F44AA1DC5E37400C9EE1B7B638E8849D23C383298E",
INIT_15 => X"015998B28654565A003F0068E35352C1CAE48BFBF3A6C9B7B286B4DA8B93D037",
INIT_16 => X"009000040A8000452110A8442040D655602A102A0027E2C42320284086E6A2EE",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"1451451E96F2FC3C34F3CF3C2AC688AA263486D3260E34C0C3A7B451B0200000",
INIT_1B => X"7A7D1E9F47A7D1E9F4D14D14D14D14D14D14D14D14D14D14D14D14D145145145",
INIT_1C => X"0007D3E9F4FA7D3E8F47A3D1E8F47A3D1E8F47A7D3E9F4FA7D3E9F4FA7D3E9F4",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"428BEF087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA0000000000000",
INIT_1F => X"80175EF0004000BA552A821FFFF8000010082A954BA00003DFEF085155400F78",
INIT_20 => X"2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BA5D2E975EFF7D568BFFFF",
INIT_21 => X"AA8015400FF84001EF0000020AA5D00154005D043FF45555540000082EAABFFA",
INIT_22 => X"F5D0415410087FD74BAAAAEBFFEF557FC00AAF7AE95555A2FBE8BEFA2843DE00",
INIT_23 => X"FF002A821FFAAD5554BA087FFFF55557BD54AAF7FBC01FFA2802ABEF557BEABE",
INIT_24 => X"4AA557BFDE10A2FBEAB45F7D56AABA082A97545F7D16ABFFFFAABFEAAFF84001",
INIT_25 => X"2092000000000000000000000000000000000000000000000FFFBE8BFF080017",
INIT_26 => X"38FD7005150438F78A2DBFF0871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC",
INIT_27 => X"0925EFF7D16ABFFE38E175EF1400000BA412E871FFE38E070280024904AA1C04",
INIT_28 => X"51420101C2EAFBD7A2FFEDB55B6A080038E3DB50555412AA8ABAAADB40092492",
INIT_29 => X"2FFE8BC7BE8E38E10A28017400E38A051FF0804050BA410A1240055003FF6D55",
INIT_2A => X"BE8A2ABD74975EDBC7550E12410087FD74AAB6AABFFC7557FC00BAE3AA9257DA",
INIT_2B => X"7F7AABAEAAF780051C70824851D7A2DB50482147FFAF554971D0492E3F1C71C7",
INIT_2C => X"00E3FFEFBD70000124AA557FFDE10A2FBEDB6DF7D16AABA08249756DF7D168BC",
INIT_2D => X"FFF552AAAAAA007BC00000000000000000000000000000000000000000000000",
INIT_2E => X"74AA0800020BA550028B550855400AAF7AEBDFEF08516AB55A2D16ABEFFFFBFD",
INIT_2F => X"A8AAAAAFFC20000000021EFF7D568BFFA2AA955FF5D04020AA002A955EFAAAA9",
INIT_30 => X"E820105D003DFEF5D51420005D2ABFF45A2FBFFF55FF84000AAAAFBC0145002A",
INIT_31 => X"7BC20BAAAAE821EFAAFBEAB55F7AAA8A00AA8417400AAAE975EF0800174BA002",
INIT_32 => X"85142010AAD157545F7AEA8B5500557DF45552A82000007BD74AAF7AEBDF455D",
INIT_33 => X"0804155FFF7D568B55FFAAAAABAFF8415545000015555A2FFC00105D7BE8B550",
INIT_34 => X"0000000000000000000AAFFFDF450804020AA557BFFE10A2FFFFFEFF7D568ABA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000400000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"5295B6957FCBE0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"6DE90201BF90102103AF158E805428249851BFB2C106592088DBF8400A5055C2",
INIT_05 => X"403DA038338041EE341036BF36812841A19B68F40A807ED9C18114956FF081DB",
INIT_06 => X"00A0E2D7D3EAFF15800100FBFB333C1CBC303163670497AFF00291B3C0E20150",
INIT_07 => X"51C581123AEE54DE8008B719E61C10BBA5DAAFA9DDA1194D51E067BB00000000",
INIT_08 => X"0320A9392083056C2270E004400091181168C4D14002A110C902481FC0B42124",
INIT_09 => X"C51DFFC40C30E5F0182D0950190C0810BE00E9A76E4C6FFBE4700000B3038067",
INIT_0A => X"F7BC81C003C001674BB55B5FBB4BB4F26A19F70027CE86F047BEF19B6D94C1C1",
INIT_0B => X"0018CFC7429F326B9E822FFC00074D5A0AB033A3F330802966F74BFF8FCFB1F1",
INIT_0C => X"3EF3D3EF3D3EF3D3EF3D3EF3D3EF9E9F79E9E00185C44B91BC1740B7605040BE",
INIT_0D => X"CFEB69FF7A5F5AFFCCA787743FE67C21800367A28FC1AAF5CF6F3D3EF3D3EF3D",
INIT_0E => X"F99FD0678B87A0003000D8D02E00000000000000040025D3C21463D6BFF252D4",
INIT_0F => X"221ABD9CA854DFDD64A67D42C0F054DFDD64667D42C063E57A8F7B4594BB02C9",
INIT_10 => X"AA504801F054DFDD64A67D42C0F054DFDD64667D42C07237DFE5865F6D2BF232",
INIT_11 => X"8EAE7F5AB50D0806A9A2E0DFFF47DEDC496DA3181A0CC71440F9FBC3EFBB5AED",
INIT_12 => X"C3FC95949AEFF556EF9C75E7DCF1EB1B6E6FCDC87CB35FC94B36AECF3A33DFE5",
INIT_13 => X"AF5B6AAAE594A4C0DBFDAD94AA669809809FEFAF4157ADB55572CA527056E9C9",
INIT_14 => X"33F32ADD543430808BABAF50E1A5EB4BAEA45A250202FE0ADD39387F92B29382",
INIT_15 => X"523E865D4B1293AB6B90BF2F0E30EDEFAFD0B3FBD72E9E90D20A003FBEBF41AE",
INIT_16 => X"02F840000BCE0B6F67B3F845E017C833F6AAC02B002A2EFF22D4073DE83FB669",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9A69A6A4624C3434C0EBAEBA21B9001804F6E62029749701020B88A7CC0C0060",
INIT_1B => X"0D46A341A0D46A341A69AEBA69A69AEBA69AEBA69A69AEBA69AEBA69A69A69A6",
INIT_1C => X"00046A351A8D46A351A8D46A351A8D46A351A8D068341A0D068341A0D068341A",
INIT_1D => X"0000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"FC00AA087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA0000000000000",
INIT_1F => X"7BE8B450051401EF087FD74AA087FFFFEFF7D168B55AAD17FFFF552EBFE00007",
INIT_20 => X"F8000010082A954BA00003DFEF085155400F78428BEFAAD168A000004020AA5D",
INIT_21 => X"0004000BA552A821FF5D00020BA552A82000552A821555D7FEAB55FF80175EFF",
INIT_22 => X"5AAD17FFFFAAFBC01EF5D0015555557BFDEBA5D2E975EFF7D568BFFFF80175EF",
INIT_23 => X"55A2D1554BAA2FBE8B55A2AE80000F7D5555555D2AAAABAAAD1420BAFFFFFDF4",
INIT_24 => X"4005D043FF45555540000082EAABFF00516AA10552E820BA007FEABEF0055555",
INIT_25 => X"AE920000000000000000000000000000000000000000000000000020AA5D0015",
INIT_26 => X"7FFEF552AB8E38087FC2092147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7",
INIT_27 => X"16AA381C0A07082497FEFB6D1451471EF007BD04920871F8FC7E3D56AB6DBEDB",
INIT_28 => X"7BEFB6DEB8E175FFE38E070280024904AA1C0438FD7005150438F78A2DBFFBED",
INIT_29 => X"7D16ABFFE38E175EF1400000BA412E871FF550A00092492A850105D2A8015541",
INIT_2A => X"AADB40092FFF5FFF6DAADF7FFD7B6F1C71EF55001756D5D7BFAEBA4920925EFF",
INIT_2B => X"2007FEDBD700515556DA2DF50492A2FFEDB55B6A080038E3DB50555412AA8ABA",
INIT_2C => X"000804050BA410A1240055003FF6D5551420101C2EAFBD7145B6AA2849248708",
INIT_2D => X"B550000175EFFFFBEAA000000000000000000000000000000000000000000000",
INIT_2E => X"AB55A2D16ABEFFFFBFDFFF552AAAAAA007BC0000557FFDFEFF7FBFFF55A2D16A",
INIT_2F => X"400AAF7AEBDFEFF7D568AAA5D2A97410007BFFFFF5551555EF087FC200008516",
INIT_30 => X"A954005D2A82155087FFFFEFAAAA975EFAAAA974AA0800020BA550028B550855",
INIT_31 => X"7FEAAAA0000021EFF7D568BFFA2AA955FF5D04020AA002A955EF5D2E80010002",
INIT_32 => X"AFBC0145002AA8AAAAAFFC2000FFD57DFFFAAFFFDF55FFD1575FF5504175EF5D",
INIT_33 => X"557FE8AAA000415410007BFFF450051555EFA2FBC0000A2FBFFF55FF84000AAA",
INIT_34 => X"00000000000000000000800174BA002E820105D003DFEF5D51420005D2ABFF45",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000CFFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"080BA868803F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"42016B0C401F58495C900A4859552A611D9A640F5903B2388004004C08A06008",
INIT_05 => X"7008000E0E508C01C28640000801133060E0032801E0202000991B708280B501",
INIT_06 => X"560000000022229A60B048048120FF040000000002C44D620F0228454C838100",
INIT_07 => X"58800A001D4033A004904087F9E3901218050018024110D6771C1F90C2856828",
INIT_08 => X"3020A82929A807B3731021400058C020000A9729400D10100420480202AC2140",
INIT_09 => X"0419002D86184A01018030430700802541420440022030041A814A0080064C1F",
INIT_0A => X"0000F0CA8428642430080438408A510185A200000045C18C0E0000A0820500B9",
INIT_0B => X"311324AA2373088479105D044A1022000001835C0C30C2E21480349D00100202",
INIT_0C => X"000C2000C2000C2000C2000C2000610006100100180A8062026000DC425C0301",
INIT_0D => X"10108003C00021002046088B5001FB3650D89844703657083080C2800C2000C2",
INIT_0E => X"007E281F840C00284A17210001060D8306C18360C1380A0260CB980840080810",
INIT_0F => X"9BBEF8E50B041029075982BF3873041029079982BF39748AA0AC800014804032",
INIT_10 => X"79BFD7F7F3041029075982BF3E73041029079982BF3F632C5F96D3C11555D5D7",
INIT_11 => X"A595405FC7F1CFEBC7586C4100A53162B47FD7E39FFEECE1598702345156AEA4",
INIT_12 => X"FE037ACFB88083A99E06271BB0CA207DFDD5920057E0B001B0EBCC79932C5F96",
INIT_13 => X"2A002DD51B6F7FC4A411D1E8D44517F14EAFE36E55150016EA8DB73E39464006",
INIT_14 => X"C30351452A13D55CFFA76E928E3891F148B30399F5FB7F28C800DFA06F5DF5CA",
INIT_15 => X"57DFEAEF1005475F1D1F608819CF0EE76E12C824ADD9089715F25FAF9DB84953",
INIT_16 => X"34041A41A0000010180C02801680460FC900052FA10DC0006DA4881C110155AC",
INIT_17 => X"60D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8",
INIT_18 => X"0D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D83",
INIT_19 => X"00000000000000000020D8360D8360D8360D8360D8360D8360D8360D8360D836",
INIT_1A => X"8A28A2891182C8A82E0820825945DF675C0770B9E11807E54587BEF8B0000000",
INIT_1B => X"2552A954AA5128944AAAA28A28A28AAAAAAA28A28A28AAAAAAA28A28A28A28A2",
INIT_1C => X"000128944A25128944A25128944A25128944A25128944A25128944A25128944A",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"57FEAA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E954000000000000000",
INIT_1F => X"D568B55080028B55002E82000087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD",
INIT_20 => X"87FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AA087FFFFFFFFFBFDF45AA",
INIT_21 => X"0051401EF087FD74AAAAFFFDF45A2D16AB55F7FFFFFFF00043DE10AA843DE000",
INIT_22 => X"00804154BA55042ABEF5D7FD75FFAAD540145AAD168A000004020AA5D7BE8B45",
INIT_23 => X"10557FD7545FF8000010082A954BA00003DFEF085155400F78428BEFAA800000",
INIT_24 => X"000552A821555D7FEAB55FF80175EF5D00020105D2A97400082E95555085168A",
INIT_25 => X"24280000000000000000000000000000000000000000000005D00020BA552A82",
INIT_26 => X"E8B550000071EFB6DF7AE921C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A9",
INIT_27 => X"FFDFC7E3F1FAF55A2DF6DB7D1C002AB7D002A82028147FFFFFFFFFBFDFC7EBF5",
INIT_28 => X"003DE28B68E38E280871F8FC7E3D56AB6DBEDB7FFEF552AB8E38087FC2092087",
INIT_29 => X"C0A07082497FEFB6D1451471EF007BD0492B6F1F8F55AADF6DB7DE3F5FAFC708",
INIT_2A => X"F78A2DBFFA28407038140410492550A2ABC7497BD25FFAADF4516DBED16AA381",
INIT_2B => X"8002E9557D1C516FA28417BD5545E38E070280024904AA1C0438FD7005150438",
INIT_2C => X"00550A00092492A850105D2A80155417BEFB6DEB8E175FF5D0E0500049209742",
INIT_2D => X"FEF552E974AA082A820AA0000000000000000000000000000000000000000000",
INIT_2E => X"DFEFF7FBFFF55A2D16AB550000175EFFFFBEAA00557FFFFFFFFFFFDFEFF7FBFF",
INIT_2F => X"AAAAA007BC0000087BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AA557FF",
INIT_30 => X"FFDFFFAAD16AB4500043DEAAFFAEAAAAA08516AB55A2D16ABEFFFFBFDFFF552A",
INIT_31 => X"FFD55EFF7D568AAA5D2A97410007BFFFFF5551555EF087FC2000FFD56AB45A2F",
INIT_32 => X"50028B550855400AAF7AEBDFEFA280154BA550400000552AA8B45087FC01EFA2",
INIT_33 => X"5D2E974000804154BA082A975EF5D517DEAA007BD5545AAAA974AA0800020BA5",
INIT_34 => X"00000000000000000005D2E80010002A954005D2A82155087FFFFEFAAAA975EF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000400000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000010228001000000000000000000024001620280000000000354200004008",
INIT_04 => X"00016200001310090090004840004152C7208802590000388000004C08006000",
INIT_05 => X"7008000E0200000000000000000100302000000000E02000009900000000B100",
INIT_06 => X"00000000000000100000000000001B040000000002C42010010200004C838100",
INIT_07 => X"E0050A040041593104004500480090080A011202201400204204018000000000",
INIT_08 => X"30E409080188000021A0000100004082A140102B4020109801A4CE0037100100",
INIT_09 => X"00000005861840000000004301000B000000000001C1C0000000000000020C01",
INIT_0A => X"0000B0C0000000101400040C0408100000000000004540800000000000000099",
INIT_0B => X"000010000800011000000000000000000000BC0007C00008092C800080000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"08000EC0000000000000000010004B2000000000000000000000000000000000",
INIT_0E => X"0006280180040000000000000000000000000000000000000000000000000001",
INIT_0F => X"4451B81A70AB3006BA0011400760AB3006BA0011400680F02096834820000000",
INIT_10 => X"04082248A0AB3006BA0011400160AB3006BA0011400084C780687DBA82800808",
INIT_11 => X"796E80A00802301BC0A7531EDD98E73B02800804620D030F873EB49F30B80112",
INIT_12 => X"0000002044F091A860700FF9198AA115D5DA37F7A80C8A3604001C0664C78068",
INIT_13 => X"51AC9000000000314E01F9F30198600631448410A2A8D64800000081B0A936B0",
INIT_14 => X"0303842281C80A23004411AD661891F15148A4420804241526D6000000000985",
INIT_15 => X"35F3D282000C6C5456C84850F61050C411AD6284FDA861682805A04A1046B2E0",
INIT_16 => X"00000000000000000000000000004600C0013800003088004202304366A4A9D3",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"86186186851046260A9A69A6039045DD1F863808633005010063A20C90000000",
INIT_1B => X"930984C26130984C261861861869A61861861861869A61861861861861861861",
INIT_1C => X"0000984C26130984C26130984C26130984C26130984C26130984C26130984D26",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"E95400F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BA0000000000000",
INIT_1F => X"FBFDFFF552E974BAA2FFFFE10087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082",
INIT_20 => X"87FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAAF7FFFFFFFFFFFFFFFFF7",
INIT_21 => X"080028B55002E82000F7FFFFFFFFFFFFDFEFA2D568B550004001EFAAAEA8ABA0",
INIT_22 => X"FF7FBE8B55AAD16ABEF5D2ABFF55080402010087FFFFFFFFFBFDF45AAD568B55",
INIT_23 => X"00AAFFFFEBA087FFFFEFF7D168B55AAD17FFFF552EBFE00007FC00AAF7FFFFFF",
INIT_24 => X"B55F7FFFFFFF00043DE10AA843DE00557FFDFEFA2D16AB55A2FFFDFEF5D2EBFE",
INIT_25 => X"04AA000000000000000000000000000000000000000000000AAFFFDF45A2D16A",
INIT_26 => X"FDFFF5D2A954AA082A92428E3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA00001",
INIT_27 => X"FFFFFFFFFFFDFEFF7F5FAFC7492A974AAB6F5F8E101C7FFFFFFFFFFFFFFFF7FB",
INIT_28 => X"00001FFBEA4A8AAA147FFFFFFFFFBFDFC7EBF5E8B550000071EFB6DF7AE92EBF",
INIT_29 => X"3F1FAF55A2DF6DB7D1C002AB7D002A82028FFFFFFFEFF7F1F8FD7AAD16AB4500",
INIT_2A => X"087FC2092F7FBF8FC7E3F5EAB45B6DF6FBEF5D2AB8F7D000000010087FFDFC7E",
INIT_2B => X"DBEF5F8FD7412ABFE28B6F5F8E820871F8FC7E3D56AB6DBEDB7FFEF552AB8E38",
INIT_2C => X"00B6F1F8F55AADF6DB7DE3F5FAFC708003DE28B68E38E284971F8FC7AAD56DB6",
INIT_2D => X"FEF552E954AA0004000AA0000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFDFEFF7FBFFFEF552E974AA082A820AAA2FFFFFFFFFFFFFFFFFFFFFD",
INIT_2F => X"175EFFFFBEAA00A2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00557FF",
INIT_30 => X"56AB45AAD56AB450004001EFFF842AAAA557FFDFEFF7FBFFF55A2D16AB550000",
INIT_31 => X"0402000087BFDF45AAD568B55AAFBFDFEF55042ABEF002A800AAF7FBFDFEFF7D",
INIT_32 => X"FFBFDFFF552AAAAAA007BC0000FFFBE8B55AAD168B55F7FFFFFFF552AA8BEF08",
INIT_33 => X"08556AB55A2D57FFFFF7D568B45002ABDEAAFFD16AA0008516AB55A2D16ABEFF",
INIT_34 => X"0000000000000000000FFD56AB45A2FFFDFFFAAD16AB4500043DEAAFFAEAAAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000800000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"0001E6000053300B00D0005800000000000000407B0004BB830004DC3D01E000",
INIT_05 => X"F0FF433EFE022001C81080001101F977E0201C409BE1F10623BB000A100CF300",
INIT_06 => X"0F00100002E22EB440012C809B2FFF7C8E8840155FDC0000010E40087D8787A1",
INIT_07 => X"3B800000000000000008407FC800B0000000100600040000C205FF91C000F800",
INIT_08 => X"28C0B0300020852000002101554021F000000000000000090492260200002000",
INIT_09 => X"00000007BEFBC010002008FF7F00000000010018A81000041C401000004FFDFF",
INIT_0A => X"0002B7C0000008000000200000200A0C004408C2007D5FC800000240001227FB",
INIT_0B => X"000000000000000000000000800800A400000000000000008000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000800080000000",
INIT_0D => X"001000000100000020000800101FFB6000000000000000000000000000000000",
INIT_0E => X"07FE29FF800C00000001002040000000000000020480002E42429C0000080000",
INIT_0F => X"4D4E180010040000400000001E60040000400000001E6010003C000000000030",
INIT_10 => X"000094B1E0040000400000001E60040000400000001E60804000000400000000",
INIT_11 => X"02000000000033628000100100000004000000006170C0008001000004000000",
INIT_12 => X"000000295810000000A100020614148002000000000004307CC3CC0000804000",
INIT_13 => X"2000000000014AC000120200000000003F0D800020100000000000A4B0020000",
INIT_14 => X"0C0C00000000002E2D000001006204040000000005786C004000000000052580",
INIT_15 => X"0A0C0939BEE1810080200000E0CE0EC000010020000000000000AE8A00002002",
INIT_16 => X"8040400400C08080000000000049F6FFC0100000000000008008008000400010",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000200",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C30C320624C1090D0F3CF3CD038001801C10000804482A60D09008269020010",
INIT_1B => X"86432190C86432190CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2C30C30C3",
INIT_1C => X"000432190C86432190C86432190C86432190C86432190C86432190C86432190C",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"4174BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA0804020100000000000000",
INIT_1F => X"FFFFFEF552E954AA000400000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA000",
INIT_20 => X"87FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFFFFFFFFFFFFFF",
INIT_21 => X"552E974BAA2FFFFE10FFFFFFFFFFFFFFFFFFFFFBFDFFF5D2E954BA007FC00BA0",
INIT_22 => X"FFFFFFFFEFF7FBFFF550800020BAAAD56AAAAF7FFFFFFFFFFFFFFFFF7FBFDFFF",
INIT_23 => X"EFA2D57DE10087FFFFFFFFFFFFFEFF7FBEAB450804001EFAAD57FEAA007FFFFF",
INIT_24 => X"FEFA2D568B550004001EFAAAEA8ABA5D7FFFFFFFFFFFDFEFF7D56AB450000021",
INIT_25 => X"5000000000000000000000000000000000000000000000000F7FFFFFFFFFFFFD",
INIT_26 => X"FFFEF552A974AA0000104AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA08000",
INIT_27 => X"FFFFFFFFFFFFFFFFFFBFDFEF5D2E974AA000A07000E3FFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974AA0071C50BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA082A92428087",
INIT_29 => X"FFFFDFEFF7F5FAFC7492A974AAB6F5F8E10E3FFFFFFFFFFFFFFEFF7FBFFFFF55",
INIT_2A => X"B6DF7AE921C7FFFFFFFFFBFDFEFE3F5F8F450004050AABEDF6FABAEBFFFFFFFF",
INIT_2B => X"7EBD168B450804021FFB6D57DE28147FFFFFFFFFBFDFC7EBF5E8B550000071EF",
INIT_2C => X"00FFFFFFFEFF7F1F8FD7AAD16AB450000001FFBEA4A8AAA497FFFFFFF7FBF8FC",
INIT_2D => X"FFF5D2A954AA0800174100000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFDFEF552E954AA0004000AAFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974AA082A820AA087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410A2FFF",
INIT_30 => X"BFDFEFFFFFFDFEF5D2E954AA0051554BA557FFFFFFFFFFFDFEFF7FBFFFEF552E",
INIT_31 => X"FFFFEBAA2FFFFFFFF7FBFDFFFFFD568B55002A954AAF7D568A00AAFFFFFFFFFF",
INIT_32 => X"2D16AB550000175EFFFFBEAA005D7FFFFEFF7FBFDFFFAAD16AB450804174AAFF",
INIT_33 => X"087BFDFEFF7FFEAB45A2D568B550804001EFF7D57DEBA557FFDFEFF7FBFFF55A",
INIT_34 => X"0000000000000000000F7FBFDFEFF7D56AB45AAD56AB450004001EFFF842AAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"1094EC681244819000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"0001E6000053300F01D4587800446194F49020107F0012BBC00202DC3823EA82",
INIT_05 => X"F0F807BFFE000120080002341881F3FFF012412A9FE1E01013BF09404050F300",
INIT_06 => X"08808210996035A000006EC2E04FFFFC0A0000101FFE4036450E08247F878703",
INIT_07 => X"003400812A156C002822987FC830F40134CC74D002016612DE87FFE004008040",
INIT_08 => X"02348D2D00080C0C53400044114000000D022640B42406808790055043A82824",
INIT_09 => X"080AC707FEFBC110008420F7FF388B70A20389346FE8000580200800008FDFFF",
INIT_0A => X"4636FFC00080013029811240444A82422A828C03BC7D7FC15025B1AB6E85A7FF",
INIT_0B => X"2019480E63180855A492712CC01C49C20201BFE45FF0C004041DA2218A8A3151",
INIT_0C => X"648A3648A3648A3648A3648A366451B2451B210018C241102068006C620C0388",
INIT_0D => X"80050094104431200090080C621FFBE0008A94641165448C80C103648A3648A3",
INIT_0E => X"9FFEADFF8050250010030165290008800440022201082401A002000C48000201",
INIT_0F => X"48A004A6C0D2820302C005A83480D1820302A009B02B101390C0CB2830816202",
INIT_10 => X"8904831400D1820302C005A83480D2820302A009B02B021A85C0941150013180",
INIT_11 => X"8834600024D052C1051E0B92D400360520202682C19024B6164E300448510140",
INIT_12 => X"4093E22A2012418A9D1D44ADD9E0F174103820101C0B8160D5516259FA1A85C0",
INIT_13 => X"8AA288209E615100280DA0052000C5006402000206C55144104D510CC1B0D640",
INIT_14 => X"D50020C04023033C52009144231D902818100C90058010361AC808126C88660D",
INIT_15 => X"2386454988140600C0181500A13E830011008B0374007000B4E0CD00024500A0",
INIT_16 => X"0224004002000000703804008001F7FFF01B982B01258088C008CC41198A1220",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"0000000000000000002008020080200802008020080200802008020080200802",
INIT_1A => X"BEFBEFBFF7FEFEFFFE79E79FFFF7CFF77FBFFEFBFF9F7E0FDF9EFEFBF0000000",
INIT_1B => X"FF7FBFDFEFF7FBFDFEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEF",
INIT_1C => X"000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0004000100000000000000",
INIT_1F => X"FFFFFFF5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080",
INIT_20 => X"7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"552E954AA000400000007FFFFFFFFFFFFFFFFFFFFFFEF552E974BA0804000AAF",
INIT_22 => X"FFFFFFFFFFFFFFFDFEF5D2E974BA002E97400007FFFFFFFFFFFFFFFFFFFFFFEF",
INIT_23 => X"AA002E974BA087FFFFFFFFFFFFFFFFFFFFDFEF5D2A974BA082E95400007FFFFF",
INIT_24 => X"FFFFFFBFDFFF5D2E954BA007FC00BA5D7FFFFFFFFFFFFFFFFFFBFDFEF5D2A954",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E954AA080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA00000",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E954BA080A000AAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA0000104AAF7F",
INIT_29 => X"FFFFFFFFFFFBFDFEF5D2E974AA000A07000007FFFFFFFFFFFFFFFFFFFFDFEF55",
INIT_2A => X"082A924281C7FFFFFFFFFFFFFFFFFFBFDFEF5D2A974BA002A95400087FFFFFFF",
INIT_2B => X"FF7FBFDFFF552E974BA0020924BA1C7FFFFFFFFFFFFFFFF7FBFDFFF5D2A954AA",
INIT_2C => X"00E3FFFFFFFFFFFFFFEFF7FBFFFFF552E974AA0071C50BA557FFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0000020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"954AA0004000AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAFFFFF",
INIT_30 => X"FFFFFFF7FBFDFEF5D2A954BA082E800AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E",
INIT_31 => X"2E97410087FFFFFFFFFFFFFEFF7FBFDFFF5D2A974AA002E95410087FFFFFFFFF",
INIT_32 => X"7FBFFFEF552E974AA082A820AA557FFFFFFFFFFFFFEFF7FBFFFFF552E954BA00",
INIT_33 => X"5D7FFFFFFFFFBFDFEFF7FFFFFEF5D2A974BA0000020AA557FFFFFFFFFFFDFEFF",
INIT_34 => X"0000000000000000000AAFFFFFFFFFFBFDFEFFFFFFDFEF5D2E954AA0051554BA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"8632CA211E4491D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"24B000808800040439245B221373581F97B0A8D1040F92000F42000047A00E58",
INIT_05 => X"0107C4410008816B105036B4180C000811E9BF2844021B1004045E4249500449",
INIT_06 => X"0111C2D50A46AE45281502E4A2200081ADA0E054402365774611E047020008E0",
INIT_07 => X"80BD5AA4BF5C91F840C1710010344DB9A808FDFF3DE0313014A2007540401804",
INIT_08 => X"EA212D6D481ADF0CE47CA21544009007A64EBD64049D028B93D9561A48F60276",
INIT_09 => X"0E48D500400015805060040080A2A0F4A82381B4000A0905A0283800AA500200",
INIT_0A => X"4E700838460402635019FBFE7FCA13520F8AAD050402204090090319A5002004",
INIT_0B => X"040F4A944B1AA313C0022AA0011C0DC0002800134000000849BCC3240A8A7151",
INIT_0C => X"70AA070AA070AA070AA070AA072550385503800500001840000C80B410014088",
INIT_0D => X"0A9CA0D458D131652A154CAC6B600085080B14004D1594832824A070AA070AA0",
INIT_0E => X"C00044000A1EC1C44140D101A54280A14050A028500A84F02842A24C594A0687",
INIT_0F => X"59E0C4E6C256690581800F1C3E82562B0581200F1C3F08145602280402080448",
INIT_10 => X"AB8581B602562B0581800F1C3E8256690581200F1C3F1238473F121000613383",
INIT_11 => X"0E1050083750B3E4275F829547008600C030374361FA2CEE046D48122C438100",
INIT_12 => X"C012A66F61154C019511628756231018500C00203E138061565160782238473F",
INIT_13 => X"AA612C0096C37B00D1724801A0009C606D1221D104553096004B61BCC1128C4C",
INIT_14 => X"41E0F0600035842E7601C2C4AC68A98810080AA825A890225189980254CDE608",
INIT_15 => X"637E00D0A1080301401C390320188321C2C0B13890105800D520AF94870B012A",
INIT_16 => X"22F110111B281A54753AA004002601001918008C10912A4440B24E8B58234A89",
INIT_17 => X"0882208822088220882208822088220882208822088220882208822088220882",
INIT_18 => X"8020080200802008020080200802008020080200802208822088220882208822",
INIT_19 => X"8000000001FFFFFFFFC802008020080200802008020080200802008020080200",
INIT_1A => X"9E79E7BFF3FEFEBEEEFBEFBEFBEFDFEF7F47F8FBEF5EB7E6CFEFBEFBE8289144",
INIT_1B => X"7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"0003F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0800000000000000000000",
INIT_1F => X"FFFFFFF5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2A954BA0004154BAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000015400F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF552A974AA0800154AAFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"AA0000174BAF7FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0004174BAFFFFFFFF",
INIT_24 => X"FFFFFFFFFFEF552E974BA0804000AAA2FFFFFFFFFFFFFFFFFFFFFFFFF552A974",
INIT_25 => X"0010000000000000000000000000000000000000000000000007FFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2A954BA000417410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080005000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF552A974BA0000174AAFFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"0000104AAE3FFFFFFFFFFFFFFFFFFFFFFFFF552A974AA0804154BAF7FFFFFFFF",
INIT_2B => X"FFFFFFFFEF552E954BA000E124BAE3FFFFFFFFFFFFFFFFFFFFFFFEF552A974AA",
INIT_2C => X"00007FFFFFFFFFFFFFFFFFFFFDFEF552E954BA080A000AAA2FFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804000100000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF552A954BA000415400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A",
INIT_31 => X"04174AAF7FFFFFFFFFFFFFFFFFFFFFFFEF552A974BA0000174BAF7FFFFFFFFFF",
INIT_32 => X"FFFFDFEF552E954AA0004000AAA2FFFFFFFFFFFFFFFFFFFFFDFEF552E974AA08",
INIT_33 => X"AAFFFFFFFFFFFFFFFFFFFBFDFEF5D2E954BA002A820BAA2FFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000087FFFFFFFFFFFFFFFF7FBFDFEF5D2A954BA082E800AA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"5886C0201A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"0005EE040057700F40D08078500000D9218020407F0000BB8018A2FC380BEAC2",
INIT_05 => X"F0F817FFFE400800020224000405F7FFE0124002FFE1E0C517FF09111212F300",
INIT_06 => X"400000409120338860900482404FFFFC000000001FFC0832050E00047F97870B",
INIT_07 => X"00246801C41C3E81E872C8FFE900FC31348EFDF03BE15E22DA07FF92C2041020",
INIT_08 => X"6220280D2B025988311AB14155421006891A1089F6E200000022C140068EB902",
INIT_09 => X"0002021FFEFBC80000000077FF184B03010004002FE1F2900201000000FFDFFF",
INIT_0A => X"0006FFEA002020626995FBE077430001E7320006F87D7FA84024B0225A890FFF",
INIT_0B => X"241C482B20400CC52492710CC80060020A81BFE41FF0C2060481200180000000",
INIT_0C => X"040430404304043040430404304021820218210018C24110A860006C620C0312",
INIT_0D => X"001002001804800000952800001FFBF040C088669070510C90C1430404304043",
INIT_0E => X"1FFEAFFF805025E00853B92588000400020001000020A8018008002000014030",
INIT_0F => X"148484054395E27E428002A4200397E07E422002A420100382FCC30832A16382",
INIT_10 => X"788417000397E07E428002A4200395E27E422002A420110A51C01C0590401486",
INIT_11 => X"1A2490040590C08120558C1759BE1C05A0400383808800DA1929F728641100C0",
INIT_12 => X"00136006000215EA0A4833A32C8832050028603050014031B3950000C90A51C0",
INIT_13 => X"658280009A2030108B14AC05C00112405222088B8332C140004D101800CE7200",
INIT_14 => X"B6808060201281004228996085F10020180C030880D11019CE4000026C00C006",
INIT_15 => X"49DC7143F01C04240030720641E0A028996483A17204680410A04104A2659196",
INIT_16 => X"1000080080000000000002001201F7FFC0011C2F81A48080CA32800A0108152A",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"0000000000000000000040100401004010040100401004010040100401004010",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974AA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E954AA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"AA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080402010FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2A954BA000015400FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E954AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080005000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA080002010FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2A954BA080407000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954BA000417410FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974AA000402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E954AA000400010FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2A954AA080017410FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2A954AA08",
INIT_33 => X"F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA080015410FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000F7FFFFFFFFFFFFFFFFFFFFFFFFF552A954BA000415400",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"0000745C200801000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"0001E6000053300F00D0007810042140C00000407F0000BB800000DC3801EA00",
INIT_05 => X"F0F8033FFE000000000000000001F17FE01240009BE1E00003BF00000000F300",
INIT_06 => X"000000009120110020100002404FFFFC000000001FFC0000010E00007F878701",
INIT_07 => X"00102050840950002802C87FC800FCAA035400001B918600C207FF8000000000",
INIT_08 => X"6234AD280B02500063AC2840001610020408178B600C24000136496087300042",
INIT_09 => X"00000007FEFBC00000000077FF000B00000000002FE0000000000000000FDFFF",
INIT_0A => X"0006FFE80000015406A800003388000025000002387D7F804024B0224A8107FF",
INIT_0B => X"20502000200000400490510CC00040020201BF441FF0C0000000000180000000",
INIT_0C => X"040030400304003040030400304001820018210018C0411020600048620C0300",
INIT_0D => X"800B00000000000000000000001FFBE0008080641060400C00C0030400304003",
INIT_0E => X"1FFEADFF80002080000000208800000000000000000020018000000000000004",
INIT_0F => X"009181008024A00043601100210024A00043C0110020901382CCCB28B0806202",
INIT_10 => X"040A03080024A00043601100210024A00043C01100209240C840C201D0210840",
INIT_11 => X"A604E0080820009908008341B000A8212070082002890010068320860C920180",
INIT_12 => X"00800082041205EC00044C1ACB66C37542082030281E0580001012811A40C840",
INIT_13 => X"27A004300004103160DB3005E000618040C022000593D002180002090166B406",
INIT_14 => X"FF20406040084210C062000C2A2DDD00180C04504086002CD680C0100010480B",
INIT_15 => X"04295C98F80400008040CC0582169022000C2876C404780028500160880012BB",
INIT_16 => X"0000000000000000000000000001F7FFC001B823018F00880008805241060208",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9EF9EFB263CC3090CABAEBAFF96857757B73E6089966B9EF9D5A220CC8000000",
INIT_1B => X"0F0783C1E0F0783C1EFBEFBEFBE79E79E79E79E79EFBEFBEFBEFBEFBEF9EF9EF",
INIT_1C => X"0000783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020100000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000400010FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2010000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA000002000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974AA000400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000400000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020100000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0002010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA000002000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA00",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000002010FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974AA000402010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00004000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"4909E6093253306F82D0007C80000000080E01007F8020BBC00040DC3801EA00",
INIT_05 => X"F0F8033FFF0240012C1400080291F17FF01241009BE1E00203BF80800000F392",
INIT_06 => X"0DC00CC0992033A062116E82404FFFFC0E0801101FFC0000010E08A07FC78701",
INIT_07 => X"00000000000000002802C87FC800F8000000000019810600C207FFF3C410D841",
INIT_08 => X"E8002000080281000008A0000014100200081000000000080480AE0000002000",
INIT_09 => X"80040007FEFBE031018C31F7FFBAEBC0020008086FE0000100280800000FDFFF",
INIT_0A => X"0006FFF800C04000000000003300800005000032387D7FE94FBEF2B2CB8DA7FF",
INIT_0B => X"20100000200000400490D10EC00040220201BF441FF0C0600000000180000000",
INIT_0C => X"04003040030400304003040030400182001821001DCCC31222730A49620C0300",
INIT_0D => X"000000000000000000012800001FFBE0008080641062400C00C0030400304003",
INIT_0E => X"1FFEADFF805025C0304001E58906088304418222C108A009A090400000000000",
INIT_0F => X"00100100000480000200100000000480000200100000100380F0C30830A06302",
INIT_10 => X"0008000000048000020010000000048000020010000000004040000010000000",
INIT_11 => X"0004000000000008080000011000000020000000020000000001200000100000",
INIT_12 => X"000000800002018C010000020800000800122000000004004000008000004040",
INIT_13 => X"2080000000040000001020020000000000800200001040000000020000021000",
INIT_14 => X"1000008001000000800200000021000020100000000200004200000000100000",
INIT_15 => X"0008400000000605000000000200000200000020400000000000002008000002",
INIT_16 => X"226410410346010000000400A011F7FFE0031823010400800000800001840000",
INIT_17 => X"2088220882208822088220882208822088220882208822088220882208822288",
INIT_18 => X"0882208822088220882208822088220882208822088220882208822088220882",
INIT_19 => X"17FFFFFFFFFFFFFFFFE088220882208822088220882208822088220882208822",
INIT_1A => X"0492410A048029890AD34D35FDD144A50CB5462D14997BE09E760AED04040000",
INIT_1B => X"6231188C46231188C49249249249249249249249241041041041041041049241",
INIT_1C => X"000B158AC562B158AC562B158AC562B158AC562B158AC562B158AC562B1588C4",
INIT_1D => X"0000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080000010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0400000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080400010FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"94A7B2B1450000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"6FEBEF5FEC737AFBC6F85FDEB220109E1FEFFFE3FBA7FDFB9BD301DC3FF5F0D2",
INIT_05 => X"F0FFEB3EFFF7FDED3FBFF6A84383F177F5FB7FF59BE1FF980BBBB7FE6D21F3DB",
INIT_06 => X"FBE564C71268F3BBF5FBFC2A427FFF7C3E3A74667FDDB7FB870FF30FFDEF87F5",
INIT_07 => X"3BC18306396FBEC14489737FDC00B13BB79DFDB83BF4112AF205FFBDD3AFB93A",
INIT_08 => X"21E4391909B381B0B1F8E041051831FA3068D77E000030021324620C0B9C2060",
INIT_09 => X"D13D980FBEFBEBF30B8D79FF7F451F33CFD60FE8FFFDF54003B1D4223B4FFDFF",
INIT_0A => X"B5AFF7CFACFAFE776F39FF7077E29D83CFAB300B017F5FFE6FBEF73BEFB967FB",
INIT_0B => X"737AF3FD62601EDC25B3533DCEB07F262213FFC67FF1C7FBFB5EC9478D5DA3A3",
INIT_0C => X"5E3035E3035E3035E3035E3035E981AF181AE315BDDCC3B336F7C548667D47B7",
INIT_0D => X"100C0E60FB9FC3A80EF69A004DFFFF7FF5F9A06E19F4DA0E80E903DE3035E303",
INIT_0E => X"7FFFF9FF8FAFAA3ADEBFB9726BAF5FD7AFEBD7F7EFFD7ACDB7F947F0EA035CF6",
INIT_0F => X"0080A40403E8BD8002000FC02003E8BD8002000FC02010979AFFE36C36B86702",
INIT_10 => X"EE00034003E8BD8002000FC02003E8BD8002000FC020037B0040A00010003E02",
INIT_11 => X"C00400003D80008160400FD81341C00020003B80008C00801EF0285380100000",
INIT_12 => X"81038406809677FA080468C46A81080581002000780C8001C8100201037B0040",
INIT_13 => X"90D162001C803411FC0024080001F80040026C0807C868B1000E401A01F11909",
INIT_14 => X"10503A00003E020042AC080CEB01228A80000F600080123E232130407080D00F",
INIT_15 => X"7520750001064180807868000110C02C080CFA0042400000F8800105B02013F8",
INIT_16 => X"FF7EFEEFF3EEC3FF7FBFFBCB7FFFFEFFE00BFF7FEBF420800EC0CBEE61F81008",
INIT_17 => X"F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F7FD",
INIT_18 => X"5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7",
INIT_19 => X"37FFFFFFFFFFFFFFFFF5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F",
INIT_1A => X"A61861BAF15EAA6AFC38E38EA3AD8ADE7A48F0B366429F434AA9FC376DAE4432",
INIT_1B => X"130984C26130984C261861861861861861861861861861861861861861869A69",
INIT_1C => X"0000984C26130984C26130984C26130984C26130984C26130984C26130984C26",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"1085B0B041000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"6FAB975B6470BAF386C87A9CB00000001FEF9F23E3A7BDE79B5101D23FB5C0C2",
INIT_05 => X"C8FFCB38FF35B44C25ADE72041A3F147F5FB7F759B91FB880BA3B6FE2921CBDB",
INIT_06 => X"B98420C71408D113956AFD0842FFFC7C3032646EFF1DB7FA868FE30EF1CE47E5",
INIT_07 => X"0041830600640C415004637FC4003021259CFDB01BF80028E001FF8251AB9D1A",
INIT_08 => X"200822020842203000082050000110023068D030000028200000008400000051",
INIT_09 => X"90A4880E3DF7E2FB0B8E717C7F411F3BC6D60B60FFDDE440018AC4AA3B0FD1FF",
INIT_0A => X"042787C5AC5ADC424B39FB6073D00D8048A31008017C1F826FFEF41FEEB027E3",
INIT_0B => X"7BEAF1C152201A4C05B7531D56B05B06A213FF863FF5D5F9FB5E8847A0702606",
INIT_0C => X"0D1030D1030D1030D1030D1030F0818688186B51BFDCC39732F3554866AD57C3",
INIT_0D => X"10080A20ED1D41880CC61A0044DFFC6EB5BCA06F18FC5A0E00F0038D1030D103",
INIT_0E => X"3FFE91FF98AEAA1AC6AC9A3A4AAD5B56ADAB56D5AFD572C597B147506203E8FC",
INIT_0F => X"0000260403C8948002000EC0000BC8948002000EC00010878AC3CB8AB8857202",
INIT_10 => X"EE0000400BC8948002000EC0000BC8948002000EC000097B0040200010003E02",
INIT_11 => X"400400003D80000070400DD81041400020003B80000410801AF0204180100000",
INIT_12 => X"010384008086378A080428C46A80080081002000780C800188000301017B0040",
INIT_13 => X"909042001C800409FC0020080001F80000007C0807484821000E400205D11101",
INIT_14 => X"10100A00003E020000BC0808EB01020280000F60000002BA222020407080102E",
INIT_15 => X"7520750000024080807868000100403C0808FA0040400000F8800001F02003F8",
INIT_16 => X"EF3AF6AF6389C2FE128971AB2DDDF8FFE0031B776BF4208006C0C92621F81000",
INIT_17 => X"D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B5",
INIT_18 => X"5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56",
INIT_19 => X"3FFFFFFFFFFFFFFFFFD5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D",
INIT_1A => X"0000001E0080397908000000A48710B4080240E543021B438A010825238B443A",
INIT_1B => X"4020100804020100800000000000000000000000000000000000000008200000",
INIT_1C => X"000A05028140A05028140A05028140A05028140A05028140A05028140A050080",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"8C2100804900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"02000100440408002408008002221000204116A280000F000001400000100010",
INIT_05 => X"00000000001265050080C000190002000000005C0000000A0000002C20600000",
INIT_06 => X"14016012000C405280200008001000011110012220009A88800009A880000000",
INIT_07 => X"0048912242288100800102000400010208000000040000082000002400814008",
INIT_08 => X"0A010040401080308400821155540001122448142491008A0049120408402210",
INIT_09 => X"04080A000000124058200408000880004440004080160C4100A8580099400000",
INIT_0A => X"4A50000080080E041000000008000C81000110010500002000000180001C8000",
INIT_0B => X"110091500020B408810000100200020408B0000020000081B2C208420ADA5353",
INIT_0C => X"5814058140581405814058140580A02C0A02C004800210C19808400500010009",
INIT_0D => X"10040860B188C0A80653020005A004039010280000800B00100040D814058140",
INIT_0E => X"600010000280000802050010660001000080004004900204020105302A000C42",
INIT_0F => X"0000A00000081480000001400000081480000001400000800C01082082210500",
INIT_10 => X"0000024000081480000001400000081480000001400000010000200000000000",
INIT_11 => X"4000000000000001400000080041400000000000000C00000010004180000000",
INIT_12 => X"0100000480802A40000000400000080081000000000000004800000000010000",
INIT_13 => X"1010420000002400040000080000000000024400000808210000001200010101",
INIT_14 => X"00100A0000000000028400004000020280000000000012002020204000009000",
INIT_15 => X"1000000000024080000000000010400400004000004000000000000510000040",
INIT_16 => X"8408420430E699AA42A1508104EA08000000810020000000044001AC20500000",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_19 => X"8000000000000000000010040100401004010040100401004010040100401004",
INIT_1A => X"20820800D41A8283AC618618EF1088160885001234B96061CCDEC4D205061170",
INIT_1B => X"6030180C06030180C08208208208208208208208208208208208208208208208",
INIT_1C => X"000B0582C160B0582C160B0582C160B0582C160B0582C160B0582C160B0580C0",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000000000000FFFFFFFFF00000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0803B2814D0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"26E1E905CC574828C4F85FC600000016004F77E2F887CDB80BC340DC07D1F000",
INIT_05 => X"F007E33E01D26CE43A92F2880B01F37011E93ED49BE01F1A03B8972E6D20F049",
INIT_06 => X"5AA06002026872BAE0B1282A005FFF001E1870223FC3BFC98101F109FC6780F1",
INIT_07 => X"3BC081023B233E804488527FDC008019968D74982C94110AF204001BC285A828",
INIT_08 => X"01E4191901A101B031F84000000831FA1028575A000110800124600C039C0020",
INIT_09 => X"C1111A0782082B50080508FF00048B124D4005C8AFF4154102914800110FFC00",
INIT_0A => X"B5AAF00A80A82C332D18ED301D229C82C7A93002017F405C409A42A9A51547F8",
INIT_0B => X"1158936D20601A98A10200308A002E240010BFC0600002AFFBE249420555A2A2",
INIT_0C => X"1A3401A3401A3401A3401A3401A9A00D1A00C000850400A11414C005005000B5",
INIT_0D => X"10080C60AB0F42A8046282000DBFFF13D059280201948B029029409A3401A340",
INIT_0E => X"6FFFF8000F8F80281A16A1504302058102C0816244B82A0CA25907D0AA015874",
INIT_0F => X"0080A40000283D80000001402000283D80000001402010901A7D694494192200",
INIT_10 => X"0000034000283D80000001402000283D80000001402002010000A00000000000",
INIT_11 => X"C000000000000081600002080341C00000000000008C00000410085380000000",
INIT_12 => X"81000006809076B2000040400001080581000000000000004810020002010000",
INIT_13 => X"1051620000003410040004080000000040026C00008828B10000001A00210909",
INIT_14 => X"00503A000000000042AC00044000228A8000000000801204212130400000D001",
INIT_15 => X"1000000001064180000000000010C02C000440000240000000000105B0001040",
INIT_16 => X"964C4A44A0C689FF3F9FFEC5D6DBFE0020096528A0B000000CC043EC60780008",
INIT_17 => X"6058160581605816058160581605816058160581605816058160581605816258",
INIT_18 => X"0581605816058160581605816058160581605816058160581605816058160581",
INIT_19 => X"17FFFFFFFFFFFFFFFFE058160581605816058160581605816058160581605816",
INIT_1A => X"AEBAEBFFF7FEFCFDF7FFFFFF5DE7CFCB773FFEFBFF3C7E1E779FFEFFF5060030",
INIT_1B => X"F7FBFDFEFF7FBFDFEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEEBAEBAEB",
INIT_1C => X"000FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEF",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"9E79E7BAF7DEBAFAFEFBEFBFFBFFDFFF7FCFF0FBFFDFF7EFDDFFFEFFE8000000",
INIT_1B => X"7F3F9FCFE7F3F9FCFE79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7",
INIT_1C => X"0003F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"1084B030000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"6DA986092050306382C05A1C900000001FAE89016387B2A38B5000D03FA1C0C2",
INIT_05 => X"C0FFC338FF008048240426200081F147F1FB7F289B81FB8003A396D20940C3DB",
INIT_06 => X"098000C51000910100006C00426FFC7C202060445F1F2572060FE82671C607E1",
INIT_07 => X"0001020400440C41C000617FC0003021259CFDB01BF00020C001FF8040009800",
INIT_08 => X"2000200008020000000820440000100220489020000020000000000000000044",
INIT_09 => X"8004800E3CF3E0B1118C31747F000B33820209206FC9E80000000000220FD1FF",
INIT_0A => X"000687C0044040424B39FB6073C0010048A20000047C1F804FBEF01BEE8027E3",
INIT_0B => X"204A608142002A440492530C401049020221BF861FF0C06C493C800580000000",
INIT_0C => X"04003040030400304003040030600182001821011DCCC31222730048620C4382",
INIT_0D => X"000802004815010008840800405FF864008880661874500E00E0030400304003",
INIT_0E => X"1FFE81FF880EA000400098200C04080204010200810020C180904240400340B4",
INIT_0F => X"0000040403C0800002000E800003C0800002000E8000100780C2C30830806202",
INIT_10 => X"EE00000003C0800002000E800003C0800002000E8000017A0040000010003E02",
INIT_11 => X"000400003D80000020400DD01000000020003B80000000801AE0200000100000",
INIT_12 => X"000384000006118A080428846A80000000002000780C800180000201017A0040",
INIT_13 => X"808000001C800001F80020000001F8000000280807404000000E400001D01000",
INIT_14 => X"10000000003E020000280808AB01000000000F600000003A020000007080000E",
INIT_15 => X"652075000000000080786800010000280808BA0040000000F8800000A02003B8",
INIT_16 => X"223010010308025410082404A015F0FFE003182701B420800280C80201A81000",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_19 => X"17FFFFFFFFFFFFFFFFC080200802008020080200802008020080200802008020",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000080040",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000F007FFFFFFFFFFFFFFFFFFFFFFF800",
INIT_1E => X"402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA0804020000000000000000",
INIT_1F => X"FFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000F",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFF",
INIT_24 => X"FFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974",
INIT_25 => X"2000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFF",
INIT_26 => X"FFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08040",
INIT_27 => X"FFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFF",
INIT_28 => X"2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFF",
INIT_29 => X"FFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D",
INIT_2A => X"080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFF",
INIT_2B => X"FFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA",
INIT_2C => X"00FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFF",
INIT_2D => X"FFF5D2E974BA0804020000000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFF",
INIT_30 => X"FFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E",
INIT_31 => X"0402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFF",
INIT_32 => X"FFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA08",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000FFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF5D2E974BA080402000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


end;