library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_plasma is
	port(clk             : in  std_logic;
        address_a       : in  std_logic_vector(31 downto 2);
        enable_a        : in  std_logic;
        wbe_a           : in  std_logic_vector(3 downto 0);
        data_write_a    : in  std_logic_vector(31 downto 0);
        data_read_a     : out std_logic_vector(31 downto 0);

        address_b       : in  std_logic_vector(31 downto 2);
        enable_b        : in  std_logic;
        wbe_b           : in  std_logic_vector(3 downto 0);
        data_write_b    : in  std_logic_vector(31 downto 0);
        data_read_b     : out std_logic_vector(31 downto 0));
end; --entity ram     

architecture ram_plasma of ram_plasma is
signal enable_a_lo       : std_logic;
signal wbe_a_lo          : std_logic_vector(3 downto 0);
signal data_write_a_lo   : std_logic_vector(31 downto 0);
signal data_read_a_lo    : std_logic_vector(31 downto 0);
signal enable_b_lo       : std_logic;
signal wbe_b_lo          : std_logic_vector(3 downto 0);
signal data_read_b_lo    : std_logic_vector(31 downto 0);
signal enable_a_hi       : std_logic;
signal wbe_a_hi          : std_logic_vector(3 downto 0);
signal data_read_a_hi   : std_logic_vector(31 downto 0);
signal enable_b_hi       : std_logic;
signal wbe_b_hi          : std_logic_vector(3 downto 0);
signal data_read_b_hi    : std_logic_vector(31 downto 0);
signal address_a_reg     : std_logic_vector(31 downto 2);
signal address_b_reg     : std_logic_vector(31 downto 2);
signal enable_a_lo_256       : std_logic;
signal wbe_a_lo_256          : std_logic_vector(3 downto 0);
signal data_write_a_lo_256   : std_logic_vector(31 downto 0);
signal data_read_a_lo_256    : std_logic_vector(31 downto 0);
signal enable_b_lo_256       : std_logic;
signal wbe_b_lo_256          : std_logic_vector(3 downto 0);
signal data_read_b_lo_256    : std_logic_vector(31 downto 0);
signal enable_a_hi_256       : std_logic;
signal wbe_a_hi_256          : std_logic_vector(3 downto 0);
signal data_read_a_hi_256   : std_logic_vector(31 downto 0);
signal enable_b_hi_256       : std_logic;
signal wbe_b_hi_256          : std_logic_vector(3 downto 0);
signal data_read_b_hi_256    : std_logic_vector(31 downto 0);
begin
process(clk)
begin
if rising_edge(clk) then
	address_a_reg <= address_a;
	address_b_reg <= address_b;
	end if;
end process;
data_read_a <= data_read_a_lo when (address_a_reg < x"0001000"&"00") else
data_read_a_hi when ((address_a_reg >= x"0001000"&"00") and (address_a_reg < x"0002000"&"00")) else 
data_read_a_lo_256 when ((address_a_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_a_hi_256 when ((address_a_reg >= x"0003000"&"00") and (address_a_reg < x"0004000"&"00"));
data_read_b <= data_read_b_lo when (address_b_reg < x"0001000"&"00") else
data_read_b_hi when ((address_b_reg >= x"0001000"&"00") and (address_b_reg < x"0002000"&"00")) else
data_read_b_lo_256 when ((address_b_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_b_hi_256 when ((address_b_reg >= x"0003000"&"00") and (address_b_reg< x"0004000"&"00"));
enable_a_lo <= enable_a when (address_a < x"0001000"&"00") else '0';
enable_b_lo <= enable_b when (address_b < x"0001000"&"00") else '0';
enable_a_hi <= enable_a when ((address_a >= x"0001000"&"00") and (address_a < x"0002000"&"00")) else '0';
enable_b_hi <= enable_b when ((address_b >= x"0001000"&"00") and (address_b < x"0002000"&"00")) else '0';
enable_a_lo_256 <= enable_a when ((address_a >= x"0002000"&"00") and (address_a < x"0003000"&"00")) else '0';
enable_b_lo_256 <= enable_b when ((address_b >= x"0002000"&"00") and (address_b < x"0003000"&"00")) else '0';
enable_a_hi_256 <= enable_a when ((address_a >= x"0003000"&"00") and (address_a < x"0004000"&"00")) else '0';
enable_b_hi_256 <= enable_b when ((address_b >= x"0003000"&"00") and (address_b < x"0004000"&"00")) else '0';
wbe_a_lo <= wbe_a when  enable_a_lo='1' else x"0";
wbe_a_hi <= wbe_a when  enable_a_hi='1' else x"0";
wbe_b_lo <= wbe_b when  enable_b_lo='1' else x"0";
wbe_b_hi <= wbe_b when  enable_b_hi='1' else x"0";
wbe_a_lo_256 <= wbe_a when  enable_a_lo_256='1' else x"0";
wbe_a_hi_256 <= wbe_a when  enable_a_hi_256='1' else x"0";
wbe_b_lo_256 <= wbe_b when  enable_b_lo_256='1' else x"0";
wbe_b_hi_256 <= wbe_b when  enable_b_hi_256='1' else x"0";



ram_bit_0_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA9918630DD2200000000000012800000040002000A106001180000000008003",
INIT_01 => X"80202100005CD2C7B4E6C1E566434955ED29B05AB311C477A91660C2B4D5208F",
INIT_02 => X"11840040D2AC24048604810082640D046B24CC461E01332121AD800087828206",
INIT_03 => X"080029800001E5202400B85242009129400A2A042000F22200808420C4108104",
INIT_04 => X"0FFF9D8F603C2128230010000300000242808041C004734430A038880239A811",
INIT_05 => X"020000002020000D274A4D200001018000080121202B00006004001212000000",
INIT_06 => X"C13448904109024705203C02E34808904139041A0823001024AC0285140000C9",
INIT_07 => X"AD0779C239A085FCE05801AA9E302EA48E692112240280820422814480043883",
INIT_08 => X"00008C001000080010000202A902E8120440D05040C204C2C131209008137028",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE0339694847C449F420A40C36848097824",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C084510228082000000000000020000000000000100004000108000000028006",
INIT_01 => X"22402100005000008490005046680400213C00142300E04080F4514BA066C00C",
INIT_02 => X"00000000000020044C00010000C28410230CC4480000024000A1800182C12400",
INIT_03 => X"00001000000000000810440001002000802880040000A2020000800004000000",
INIT_04 => X"006D858F60240028030010000140042911000040000032800000194004190008",
INIT_05 => X"A400000020200008014002200009080109000484820B00000000004848400000",
INIT_06 => X"010448504104201100008100002905400211220002A480048118000054040008",
INIT_07 => X"024205F019200280860000100002101406492022102200040000821212481910",
INIT_08 => X"080004204840000000080A08000A2A454002080000090A458294C24001820004",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE0614546024C1E10064251C088C4057AA0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0C0400000682101010101000092D555550554161001447421116AAAAA820012",
INIT_01 => X"0A001DAAA04408028418019800610454A10E00C4000CA262012000C8A0780028",
INIT_02 => X"100400120DC92A5D0C4335282951264102C1C140091444504A900282D2604003",
INIT_03 => X"82921220A28080400A92560001002012E062020401AE088010808000E4110B00",
INIT_04 => X"8000400010008001800040A2216AA439410080C0150120A80412106024900048",
INIT_05 => X"25280502622420C2000400A080C908191E12C4ACB24801600AA8284ACB6C0208",
INIT_06 => X"148401F4350564088D5442812C85210C221008A80880840DE318001020869400",
INIT_07 => X"025294C0908082810984424022C89D102421207614640008B4088012B2221060",
INIT_08 => X"4B3D0D0149D2C586804809008008A21544460200150B9A8D46B4AE500242A910",
INIT_09 => X"0000000000000000001FFFFFFFFFFFF62A53D68064DC5B30EAD404FCF071D0A1",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C081002008E009100110011024C366666619989C00210D460141B33333020006",
INIT_01 => X"0004B52CA4642830841112880080922C210C4480004812E055808C413181DC4C",
INIT_02 => X"101400182DD13AA94549640B18C2C44822849440480EA8148220888292050048",
INIT_03 => X"3183106A69989A5449B054A8102C240814A02200102C08101280808005100940",
INIT_04 => X"00000000104000410400408289599019410A02020D802098421090509410426A",
INIT_05 => X"E02873200000280081010000A00818001C0204ACA6C343038663254A4ACA200A",
INIT_06 => X"040C015D38052540005005141C14210422140822A0A429850A09B00002131800",
INIT_07 => X"0210048010000082068A043000C2811004010080142004006145001292801040",
INIT_08 => X"D19486014BD283038520180021088AD1514649018C298A8542BCAA5085880C80",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE450C1460054143016A2C000887031D238",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C48B20BC128580000111100000FC78787806181810000D18095E3C3C3C028006",
INIT_01 => X"0800252A604408128400100081842028A108042040C20260028008C0D0001E0C",
INIT_02 => X"920406120DD124110D42040879D2002022409100095E641048102008D2214003",
INIT_03 => X"87840669E7D0108253B6470800292C1018000000002E28001080601083130802",
INIT_04 => X"A00060000000000184010202A1B86529085010103E41203A0E02503474900026",
INIT_05 => X"60088F0A2A04610881110089810A09085C00048C828243571E19014848F0008A",
INIT_06 => X"1484017E820421508016840008A0A449401010C9832ADD24801B2400040C2100",
INIT_07 => X"0012848090001023048A4420008A9510240104A010202005E11C0612126A1010",
INIT_08 => X"DB9507014DC282878CE88108103AAE30F30E2B243C299A0D069C8E4085020880",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE949202102283E622408110054C4451803",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"CEC8381F030781111000000000D7807F8048181E94284D60B555C03FC0120006",
INIT_01 => X"082025836054C8D69416D281E46C6D2DA50DA4A0F217E665A82460C8448012AC",
INIT_02 => X"918425005D45A411060604228642890040A491061E213031012C8000D7030206",
INIT_03 => X"6860699410016D322440A8D20600910304200004210010AA4082501400108001",
INIT_04 => X"AFFF9D8F603C2169A70150280207E432004880C5C0147145B1A0788B0638B911",
INIT_05 => X"C102609A62E44401230244A910230049482021090431009161FD24109000000A",
INIT_06 => X"C1BD40D46D080351A5B0A506EB684DD140BD0611E8998218802C8012C10401E9",
INIT_07 => X"A7056C8238820158E6980032BEB03FF08E21A02A2084008A18A3860404CD3890",
INIT_08 => X"2D89A40010321280520C894819004C070000C0B34342A4120901008001817B0A",
INIT_09 => X"0000000000000000005FFFFFFFFFFFEF7800000EF9FA8F76FC3ED7FDBCFDE954",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08C0708E06000000000000000D7FF80000FE01E94A845609155FFC000100002",
INIT_01 => X"081425AC41440812842012C018610038A10804B00C14A062001000C08000100C",
INIT_02 => X"120420020080A411054204280152000008809101410220044820000080210142",
INIT_03 => X"400010080000081208585489802024C014200004012E08805082000000121000",
INIT_04 => X"0000605096408404000A00000040142940480000000020810000104204100108",
INIT_05 => X"210A401822E44400980130A91038094040202CACA6804012000065CACAFA2240",
INIT_06 => X"040D0094000521402410040008082000481400034AE2420CA009801281040000",
INIT_07 => X"401004801002102384824420008081500401A48814A4200801010432B2801000",
INIT_08 => X"09802701C9F2130806EC804230180201000A03240039AA954AB4AA5085000B82",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE83BF7F7867CEE7F72EAD507FCFC7CF8A0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4CC031862648000000000000000000000000000840844008100000000100006",
INIT_01 => X"0804250020440802842102C012099610A10040B009001060000008C014000C2C",
INIT_02 => X"10040010008024110402040001D2040000809100410220144820000090210042",
INIT_03 => X"40001008001210084840108880600C4034200000000000098080000000100000",
INIT_04 => X"0000002080004802008608000140110048080000000228810004144205140428",
INIT_05 => X"4040401020E120828905102480A310501C10A02820C040020000000202000000",
INIT_06 => X"240D23F991019008240444040088200140148002A20082088008800000040026",
INIT_07 => X"00100481140A8081848A4220200884504503A06E068400280100800080009420",
INIT_08 => X"0264260101B1D102040428480810841500040002000030D86C382C1001000312",
INIT_09 => X"0000000000000000001FFFFFFFFFFFF200000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"D4C80010020C811111111111000000000000000000800C000100000000000002",
INIT_01 => X"0804258021440812842112C000099638A10844B000141062000009C814800C2C",
INIT_02 => X"100400100000A411040204200042000000801100400220140020000090010042",
INIT_03 => X"5000000808020A1000584481840028C204200004012E0888D080000000301000",
INIT_04 => X"A000621010418645C45946AAA800100900480002000004014000020204024000",
INIT_05 => X"210A400022240000190030A80019280048000C8C9210040280002DC84DFC22CA",
INIT_06 => X"00001050032460500004840000A8044040004009000002048008801281040024",
INIT_07 => X"0000048002000000848800202008001000810026506200040101963236C80210",
INIT_08 => X"141D0401CA5011080400000210180E010006400200191A0D068C864421000000",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE74B67630200DA6122CCA8C0FCFC7D6140",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100204811111111111000000000000000084084C008100000000100002",
INIT_01 => X"0010250AA0440812840112C000609228A10044B00000B060000008C014000C2C",
INIT_02 => X"B2042780008024110402040001D2046008C00001010264104A30200292214103",
INIT_03 => X"5000100808000A100850448800202C0014200004012E088050827814C2B20003",
INIT_04 => X"A000600010408441840142AAA840100900480002000102814002414204814008",
INIT_05 => X"A10A401822C440008001008900292840480024849280441280006D484DFC22CA",
INIT_06 => X"140908D0012420502404840400A825400004208848080204A0088012C1040000",
INIT_07 => X"021084808162102084880020200884502059842A50A420480100961212CA0110",
INIT_08 => X"0000260049E010000404804030080A00200A402200092A158A94CA4421000302",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE4234A4E04D5408102225FC4FD58D98220",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100264811111111111000000000000000084884C008100000000100002",
INIT_01 => X"0810250360440812840112C000609228A10044B00000B060000808C014000C2C",
INIT_02 => X"10040000000024110402040001520000008011010102201048200000D0210102",
INIT_03 => X"4000000800000810004800880020041014200000052C00805080000000100000",
INIT_04 => X"A000600010408441840142AAA800143000480000000100010002000204800000",
INIT_05 => X"C10A401222E40000810100A8003210484800280814C0400200002D8081BE224A",
INIT_06 => X"1489005002004010A0008404002025500804000808000208A0088052C1040000",
INIT_07 => X"4210008080020001048A4020200080402001800C00C400480101062024CA0010",
INIT_08 => X"0000260081B00080040401423010040100040002001030180C180C0001000302",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE771F0778E5016F81494EC15A01C5DA140",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C2880203B0600020202020200000000000400000000004001100000000000006",
INIT_01 => X"082425AC40448882840602C168004100A10180B0B4004064000000C00000000C",
INIT_02 => X"110400121014A411074204280042010000801104540220240024000080010042",
INIT_03 => X"40000888000041002040009302000181042000000000000A8080000000100000",
INIT_04 => X"0355134A4410692C60861400000010000008000080000B0100800582072A2001",
INIT_05 => X"0000400020000000320064000000000008000000000000022000000000000000",
INIT_06 => X"802050500000000100000400420000000029400000010200802D8000000400AC",
INIT_07 => X"8C0518832A800212449004200C200A20CA81008000000000010000000004AA00",
INIT_08 => X"0004050000000000040008080800801400000012002000000000000085030080",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE7394D4E04C1148010440605A158D94040",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C88A1F83F000020022002200020000000040004000000480012A000000000002",
INIT_01 => X"081025A00054C8C6940202C06F000801A50080B037810465AA0C60C00000008C",
INIT_02 => X"110400125014A4110746042880428100008411010603302100248000C0030106",
INIT_03 => X"4000018800010400044000DB822095C1142000002000102B8080000000100000",
INIT_04 => X"0F9B1B4E8208012E62940800020010000008808100000A4120000502072F8000",
INIT_05 => X"0040400260000001BA0374000000000808000000002100024000000000000000",
INIT_06 => X"81A078504000000180002502604008800029E01000000210802D8000000400EF",
INIT_07 => X"000400832F6000410692403298002000CBD90000000000A0012200000004AF80",
INIT_08 => X"0004070000001180040001000000000000000002400000000000000001806000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE701B2B18095005C029A93123518991024",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C6CC00100206811133331111580000000000010084084480A320000000100002",
INIT_01 => X"083425A020C40812840552811060DB28A10144A08801F060003809C014000C2C",
INIT_02 => X"114400321014A4110742042803520800408011054102201449240000D4210342",
INIT_03 => X"4800000800016D300048A0880020041014200001832C10A85080020000104400",
INIT_04 => X"ACE2ED56765C846DC75B56AAAA00109204480849C007540130A62A020480A800",
INIT_05 => X"410A401226C400218203048800321448480029091490400A60042D9091BE225A",
INIT_06 => X"7599005002184000A1002402434028800004001004000208800D8032810400E0",
INIT_07 => X"A515688080020959648240201830A2E02001820C20C4104A01030C2424820080",
INIT_08 => X"0004270091B0008034044140101044020004801A0052341A8D194C821101530A",
INIT_09 => X"0000000000000000005FFFFFFFFFFFF83800001EF9FE0F76FC3ED7DDE4E5F8C0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C088000001600222000000005A0000000040014000000480012A000000000002",
INIT_01 => X"08002500004408028400828000600000A10020A00000A060000000C00000000C",
INIT_02 => X"1084000000002411040204000042000000801100000220000028000081010002",
INIT_03 => X"4000000800000000004000800000000004200000000000000080000000108000",
INIT_04 => X"000D873106394000021014000200100000080000000000010000000204000000",
INIT_05 => X"0000400020000000000000000000000000000000000000020000000000000000",
INIT_06 => X"0000001000000000000004008000000000000000000002008008800000040000",
INIT_07 => X"0000008000000000048000200600000000010000000000000100000000000000",
INIT_08 => X"0000440000000000040000000000000000000002000000000000000001000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE07BF7F78E54CEFD36FAFD17FCFC7CF320",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08800000060022222222222000000000040000000000400010A000000000002",
INIT_01 => X"08002500004408028400028000000000A10000A000000060000800C00000000C",
INIT_02 => X"1004000000002411040204000042000000A01102160220000020000080010002",
INIT_03 => X"4000298800000000244008800000000004200000000000000080000000100000",
INIT_04 => X"0000008000042B24218800000200100000080000000001450000008A04000011",
INIT_05 => X"0000400020000000000000000000000000000000001000020000000000000000",
INIT_06 => X"0000001000000200002004000000000000000400000102008008800000040000",
INIT_07 => X"0000008000800000048000200000080000210000000000020100000000000000",
INIT_08 => X"0000040000001000040000000000000000000002000000000000000001000000",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"05104816EA00C199999999998B82D55555055577C0000675C3816AAAAAB80003",
INIT_01 => X"8014102000081213688B1862C400120ADA22C61962221218A90010E0957F0E0E",
INIT_02 => X"C200BAC50001061C8901300A2C0980A50085C801003641100400A00980206443",
INIT_03 => X"E2D5423CB284889002E20281C02900E8CC00000340A9401040162E6680824001",
INIT_04 => X"DAC651494D654F010FCA0208282AB2000D98181C14FDFC29876BFE33310017A2",
INIT_05 => X"0162E5846A0444221C5838881100401021048000000145D30AA9290000198B2F",
INIT_06 => X"84140A00A840000022800281241080040000104000002F219092A594094A9406",
INIT_07 => X"00000001010104011A42801D0244100440014000800490D0B58C444000A08004",
INIT_08 => X"612A8AB000AC00B4C66130400020000011002743150000000000100000548522",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE0334A4A0C60F6FB363875D4C538399B91",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4F74BF57E6E587FFFFFFFFFF92D71999998E665DC000E1D9E8758CCCCCF80000",
INIT_01 => X"2ADE30F033C915094A13393EDEF4B2265284CE4B6F40B85001AE0AB1FA003513",
INIT_02 => X"664123B786736A3991E3A47C1D59727F83855D59A1AC21CA6C30AAA2F8F149E3",
INIT_03 => X"01EF407061DE98DF4182021FC45117E22A0888D2C6F8E0FE6823B275CDE77725",
INIT_04 => X"D90A855E9396159B5AEBFD777C19EBC03DF139380EEDFC180363FE101FCE17A2",
INIT_05 => X"078D83F7F3CEFAFFFC5FFB96EBC021EE7D7ED00008BD6BB0067A7300009CCDED",
INIT_06 => X"5FEBF17BF430142FF1415AD12C11700001FFC007E7FAE8210DCA47FF1E58E6B8",
INIT_07 => X"105801B3FEE93C0112E1DACF82C6D945FFBB0E504085A1D076041DC000A6CE27",
INIT_08 => X"E66D1FC40024DFE9C023F3F007600088771815600D0020100800010630ECAF77",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE00C363180DDE2F82193AAC100343592A0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"80900040060040000000000040039E1E1E0F80060E1C067E2F81CF0F0F000003",
INIT_01 => X"82500F0000100211A6110064200002886984501A10005048A99041D0557F0A28",
INIT_02 => X"C0404B0000108804C04211220424A28000C0804940226454001080009001A502",
INIT_03 => X"6078001C3080000000EB02801129001CDC40000100810011D008380302004002",
INIT_04 => X"A662F955E7094500A5D54008A007F014021880C4040200098204001310000002",
INIT_05 => X"5062E0880ED505001C0038001036D20000002A1A1500108301F98CA1A12F1240",
INIT_06 => X"A4150A040AC0C8020A920A081014C00C2080386000000B2A5882A400218B3806",
INIT_07 => X"00500000008200051B06814AC10000000020810D82484020198561286D113146",
INIT_08 => X"266BAC10A190201046240000001405208005018303969048A41A4C084AD08000",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE00917109AA06CA940889D014484C5D990",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"00014020080007FFFFFFFFFF82D7E01FE008005FC000E7E1C1F5F00FF0380003",
INIT_01 => X"0000000000000004108800000000000104220004006A80000000000000000000",
INIT_02 => X"00009440000005400C0000020400000000000000002200000020000940000000",
INIT_03 => X"6040001C3080000000E20280000900000C000000000000000014440010000010",
INIT_04 => X"018F03201F7C056400DE0C82A800700000180004040000098200001310000002",
INIT_05 => X"0000E08000000000000000000000000000000000000000830018000000302240",
INIT_06 => X"000000000000000000000100000000000000000000000B20831BA40000240100",
INIT_07 => X"0000000000000000000000100000000000000000000000001184000000000000",
INIT_08 => X"2110402000000000462000000000000000000103010000000000000000000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE02EDADE84C87AAA0501480081CC8CB890",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"00000000000007FFFFFFFFFF82D7FFE0000FF85FC000E7E1C1F5FFF000380003",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000027C00000180004400007E00000000000000000000",
INIT_03 => X"E7C6867DF780000093E60380000900000C000000000000000000000000000000",
INIT_04 => X"A01182938901EA66400042A800BFF000001800043F10023B8E18013770310046",
INIT_05 => X"0000EF8000000000000000090000043020040000000007CF1FF800000401401A",
INIT_06 => X"000000000000000000000000000000000000000000001F200002A40000000000",
INIT_07 => X"00000004012900000000000000001004004B400000101001F99C000000000000",
INIT_08 => X"E0040100040C4805EEE00000000000000000230F3F0000000000112000000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE0402621121D803000120200200848E033",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4410801502168D555555555520D7FFFFFF90001F8000057F8D55FFFFFFF00002",
INIT_01 => X"8880BE000439376128C090A2E09240284A30242970600098540084F0017FA04B",
INIT_02 => X"0511481A600817F8800B64437D11428202208800047EF900C80488000085480F",
INIT_03 => X"E7D80EFFF7CC20E513E60BF2044D11000C800040108C0022022B789ECAA60068",
INIT_04 => X"A339708A60102128A000100000BFF000281B33343C01007B8E02003FFA280436",
INIT_05 => X"0400FF909010C50924424A0A4E0001004202001000202BC71FF8010000B8224A",
INIT_06 => X"803440026C000403008142D00504C00C20E91842A2A29FA1D882B4013A0BC088",
INIT_07 => X"21004806380200410AC4DA18814000418A00800040002047F9DC000040152848",
INIT_08 => X"F7F9E20001A3C285CFE02200024000A2D500B307BF0020100800000000F05610",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE038888C1EF9FE0FF6FC3CD7FDFCFD78DB",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"6CD0E84501520D555555555524FFFFFFFF90009F8001C17F8055FFFFFFF00000",
INIT_01 => X"0A94BEAFE77D3C314A43D337A45241685290F4CFD22090F85C488C03D57FAC62",
INIT_02 => X"F6157F9A78589FFDD14B756901537001E028C4415900AB14E83DA22A50A5694B",
INIT_03 => X"0827A802001090086000807A1124150890A222023DA002AA52AE78DFEAF6314B",
INIT_04 => X"AFBB390A30488569A60142AAAA0003022943B3B043B10100111A80008AA81AC0",
INIT_05 => X"052A101242D56D8BA4574A886E20405943422101103308000007AC10111C264A",
INIT_06 => X"95B9400000680303A0700FD92A012001036D0602A2A68081D98111502ADFFEA8",
INIT_07 => X"84170066A882B0892642407D02A2B185AA202C00A20445CC006054040096280A",
INIT_08 => X"17FD23001023D3900105A3409342604044500400800084422111088C6164DF12",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE07B77739EF5EEFB76BAFF15E4BCFDF3A8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"8A99D0720284A800000000006A000000005FFF400C1804002D00000000000002",
INIT_01 => X"A00080000420E3E7BC8241B640909201EF20906F206006E5F4E2B4F0200040CD",
INIT_02 => X"A39050087D451C8190084003FC04B16802C11910167EDC8180382AA20006800C",
INIT_03 => X"E7C02FFFF780000017EE0BA0044D00122CC888D0700CC010020D0094F2A38B73",
INIT_04 => X"0CCAAD86201C00280300100000BFF010001A02043C0C517F8E6028BFF0000017",
INIT_05 => X"4000FFC89801B282044400068092100014108808048043C71FFF818080920000",
INIT_06 => X"41040000420040000B034B10850100000010002000013FA88082B4013ADFFF40",
INIT_07 => X"000000000008000109A00A58044208000002004400420003FDFD002024201006",
INIT_08 => X"E000800080100005CFE00000001004A091043B97FF1200000008000002F83400",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE00000000000000000000000000000001B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010800820001080000840037C00000000000000007E88008380000000040008",
INIT_03 => X"E7C0067FF780000013E603A0000D00000C800000100000000210008001000040",
INIT_04 => X"0065E581003800000200100000BFF000001A02043C00003B8E000037F0000006",
INIT_05 => X"0000FF8000000000000000000000000000000000000003C71FFF800000300000",
INIT_06 => X"000000000000000000000000000000000000000000001FA00262B40281000000",
INIT_07 => X"000000000000000000000002400000000000000000000001F9DC000000000000",
INIT_08 => X"E000400000000005CFE000000000002091002307BF0000000000000000000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE01D1A18B4B598CC60523ACB39BEBD603B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010000820001080000840037C00028600040000007E88008000000000040008",
INIT_03 => X"E7D8067FF7DC38FD53E623A0000D00000C800000100000000200008000000040",
INIT_04 => X"0000600C600421202100000000BFF000001A02043C00203B8E001037F0100426",
INIT_05 => X"0000FF8000000000000000191120214040200010000027D71FFF890105B40080",
INIT_06 => X"0000032FBC009428008000005014C00C2080184000001FA00002B40000000000",
INIT_07 => X"A5414910100200586004900081100AE00400800840802001F9DC000040010060",
INIT_08 => X"E002201C05A0000DCFE00000002000229108A327BF0230180C100C0000002200",
INIT_09 => X"0000000000000000003FFFFFFFFFFFE020272920E9ED0B200C52CF20B83A81DB",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"85F820440E61E5DDDDDDDDDD81D7FFFFFF8FFE3FDEBCEF7FDFD5FFFFFFF80007",
INIT_01 => X"AA5E3FF033CC1A1BA4993AAC8064328EE9265EAA400ABA7000401AC1DE00573E",
INIT_02 => X"F645FFF78F73EF7DDDE3B57E7C6F72BF89C15D49E0FE675E24302AA9F8D1E5E3",
INIT_03 => X"E7FFD67DF7DE1ADFDBEF578C5479263E7E600053CEFDE25C78BFFE7FDFF77F3F",
INIT_04 => X"F000600019C294D19C21E3FFFDFFFBDD7FF9393C3FF980BB8F5BC0777CC057EE",
INIT_05 => X"76AFEFFFBFDFFFFEC44D899FFFFFFFFE7D7EFEBEBFDE7FFF1FFBFFEBEFFFFFFF",
INIT_06 => X"1ECB83FFBFF5FD6EFED75ED91C9CF11D68861AE7475A7F2FDFDBE7EFBFFFFF30",
INIT_07 => X"525A85B4C00BBCA59DE7DBED41CEC5553003EF7FD6FFF159FF9DFDFAFFB34067",
INIT_08 => X"FFFFFFFDEFFFFFFFEEEFF3F2377C0F29F31F676F3F9DBA9D6EAEBF7E7B7C8F77",
INIT_09 => X"0000000000000000003FFFFFFFFFFFE0034B422CD53444E373420BBD2C2CFAB3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"11200008002844CCCCCCCCCC80D7FFFFFF8FFE1F5AB4AB7F5ED5FFFFFFEA8015",
INIT_01 => X"080A0E5012800008002029000029049200080A4000142822000002090A800110",
INIT_02 => X"4441D8370DC3416110A004547C8854AB88011100A0FC000A040022202A1000A0",
INIT_03 => X"97EF9671EFDC1ADDDB97570404512A062A000057CA7F0844783D024B19456E38",
INIT_04 => X"F000600019C294D19C21E3FFFDFFEEED6471292A3FB880BA4F598074784056EE",
INIT_05 => X"B08F8FF597FFB2B2410480BECEADCE767554B6B6BBCC7BEC9FFBBF6B6BFDFF7F",
INIT_06 => X"0E4383AFBDD5BD7A76D7C05C1CACF55C688218EC0C023C267842452AEBF3DE10",
INIT_07 => X"5A189424400B2A2290A9DE0561CCC5511002CAEB96BD5119FE1CEE9ADBF94076",
INIT_08 => X"FFFF31FD6BEFE677E8EF78FA3E4C8B1D1113474C3F2DAA956AA6BB7AD42E0FD3",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE03F1110E441278421012A097022228883",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4128400000606088888888888000000000000000420526004380000000080003",
INIT_01 => X"220A20501184080808802A90006000C202200AA40000A820004A02822A004110",
INIT_02 => X"B24427A5000A440440A21114001A00002288C440A980220A0CA1088828B120A2",
INIT_03 => X"0000000000008000800100041110020C8222220186D182D428827A14E2B25403",
INIT_04 => X"50000000098210901820A155540009C40D2018180000A0000001100000500000",
INIT_05 => X"15A5002D0D0A4D38405082013104A72722261202091E1438000012202401D9B5",
INIT_06 => X"0A46800000B00800500004000001100103520206A6A480028100406810240010",
INIT_07 => X"104A014050019880140100200006500414006601401B30140200388809005000",
INIT_08 => X"0000D0E0240C34682002D2B0852621C8444918E8000400400012112631000041",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE02064636888C821822C1405C480005B40",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A5F0A0540E75C5DDDDDDDDDD81000000000FFE20C60C677EC3D5FFFFFFD80003",
INIT_01 => X"805E1FFFF1C81619E659392E8076B2AE79965E4B402AB858000A0A71FF7FBF3B",
INIT_02 => X"E240FFF78F72EB588DE1A03E016D627D81408809E0FE455E66100001F850C5E1",
INIT_03 => X"E037C67C104E00C793E9038C403806345E4000438F5D604C281FFE7FDFA35F3F",
INIT_04 => X"F0000000098210901820A15554BFFBD43EB9191C03F1A03B811BD0370CD013C6",
INIT_05 => X"5285E07FAFDEDDF4C409891B75D6B6EE3D3C5A0A0D9C1FFF0003F2A0A4BFFBFF",
INIT_06 => X"1ACE817992B0592EDA015AC90010100001160005455A5F0B5E9BE3FFAE2BE130",
INIT_07 => X"100800B0D0011C0519C74BCC4004400034014755405DB059FF813DE82D92502F",
INIT_08 => X"17FFDFE8A4BFFFEDEE03D1B0173405A8A20D37EF00941008040A15263A748175",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE0F480845EF1DE1EFDF8B9DEFDFCFDF890",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000222222222225A00000000000140000000800020000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE03B7F7BFCFDFCEFE37F7E0FFDBCBDF3E0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"60008010001404444444444400D7FFFFFF8FFE1F0810817F0C55FFFFFFE00000",
INIT_01 => X"08800E0FC20105004A40000200128020129000010020000800000030017FA801",
INIT_02 => X"4401D8120D410161100004407D1050EB80011110017C00804A00222200200800",
INIT_03 => X"87EF8671E7DC18DD5386030004410002280888D2492C0080503D004B19452A38",
INIT_04 => X"A000600010408441840142AAA8BFE200205121203FB8003A0F588034780016E6",
INIT_05 => X"010A8FD092D5B2820004009ECEA040505450A01010806BC41FFBAD0101BC264A",
INIT_06 => X"0401032FBC40952822D340581C04E00C20C0186000003C2058420512ABD3DE00",
INIT_07 => X"00100004000A200000A0DA0541C081410002884882844109F81C440040B1006C",
INIT_08 => X"F7FF211C01A3C215C8E5204012400000111007043F00A05028100808402C0F12",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE000000000000000000000000000000003",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA9918630DD2200000000000012800000040002000A106001180000000008003",
INIT_01 => X"80202100005CD2C7B4E6C1E566434955ED29B05AB311C477A91660C2B4D5208F",
INIT_02 => X"11840040D2AC24048604810082640D046B24CC461E01332121AD800087828206",
INIT_03 => X"080029800001E5202400B85242009129400A2A042000F22200808420C4108104",
INIT_04 => X"0FFF9D8F603C2128230010000300000242808041C004734430A038880239A811",
INIT_05 => X"020000002020000D274A4D200001018000080121202B00006004001212000000",
INIT_06 => X"C13448904109024705203C02E34808904139041A0823001024AC0285140000C9",
INIT_07 => X"AD0779C239A085FCE05801AA9E302EA48E692112240280820422814480043883",
INIT_08 => X"00008C001000080010000202A902E8120440D05040C204C2C131209008137028",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE0339694847C449F420A40C36848097824",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C084510228082000000000000020000000000000100004000108000000028006",
INIT_01 => X"22402100005000008490005046680400213C00142300E04080F4514BA066C00C",
INIT_02 => X"00000000000020044C00010000C28410230CC4480000024000A1800182C12400",
INIT_03 => X"00001000000000000810440001002000802880040000A2020000800004000000",
INIT_04 => X"006D858F60240028030010000140042911000040000032800000194004190008",
INIT_05 => X"A400000020200008014002200009080109000484820B00000000004848400000",
INIT_06 => X"010448504104201100008100002905400211220002A480048118000054040008",
INIT_07 => X"024205F019200280860000100002101406492022102200040000821212481910",
INIT_08 => X"080004204840000000080A08000A2A454002080000090A458294C24001820004",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE0614546024C1E10064251C088C4057AA0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0C0400000682101010101000092D555550554161001447421116AAAAA820012",
INIT_01 => X"0A001DAAA04408028418019800610454A10E00C4000CA262012000C8A0780028",
INIT_02 => X"100400120DC92A5D0C4335282951264102C1C140091444504A900282D2604003",
INIT_03 => X"82921220A28080400A92560001002012E062020401AE088010808000E4110B00",
INIT_04 => X"8000400010008001800040A2216AA439410080C0150120A80412106024900048",
INIT_05 => X"25280502622420C2000400A080C908191E12C4ACB24801600AA8284ACB6C0208",
INIT_06 => X"148401F4350564088D5442812C85210C221008A80880840DE318001020869400",
INIT_07 => X"025294C0908082810984424022C89D102421207614640008B4088012B2221060",
INIT_08 => X"4B3D0D0149D2C586804809008008A21544460200150B9A8D46B4AE500242A910",
INIT_09 => X"0000000000000000001FFFFFFFFFFFF62A53D68064DC5B30EAD404FCF071D0A1",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C081002008E009100110011024C366666619989C00210D460141B33333020006",
INIT_01 => X"0004B52CA4642830841112880080922C210C4480004812E055808C413181DC4C",
INIT_02 => X"101400182DD13AA94549640B18C2C44822849440480EA8148220888292050048",
INIT_03 => X"3183106A69989A5449B054A8102C240814A02200102C08101280808005100940",
INIT_04 => X"00000000104000410400408289599019410A02020D802098421090509410426A",
INIT_05 => X"E02873200000280081010000A00818001C0204ACA6C343038663254A4ACA200A",
INIT_06 => X"040C015D38052540005005141C14210422140822A0A429850A09B00002131800",
INIT_07 => X"0210048010000082068A043000C2811004010080142004006145001292801040",
INIT_08 => X"D19486014BD283038520180021088AD1514649018C298A8542BCAA5085880C80",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE450C1460054143016A2C000887031D238",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C48B20BC128580000111100000FC78787806181810000D18095E3C3C3C028006",
INIT_01 => X"0800252A604408128400100081842028A108042040C20260028008C0D0001E0C",
INIT_02 => X"920406120DD124110D42040879D2002022409100095E641048102008D2214003",
INIT_03 => X"87840669E7D0108253B6470800292C1018000000002E28001080601083130802",
INIT_04 => X"A00060000000000184010202A1B86529085010103E41203A0E02503474900026",
INIT_05 => X"60088F0A2A04610881110089810A09085C00048C828243571E19014848F0008A",
INIT_06 => X"1484017E820421508016840008A0A449401010C9832ADD24801B2400040C2100",
INIT_07 => X"0012848090001023048A4420008A9510240104A010202005E11C0612126A1010",
INIT_08 => X"DB9507014DC282878CE88108103AAE30F30E2B243C299A0D069C8E4085020880",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE949202102283E622408110054C4451803",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"CEC8381F030781111000000000D7807F8048181E94284D60B555C03FC0120006",
INIT_01 => X"082025836054C8D69416D281E46C6D2DA50DA4A0F217E665A82460C8448012AC",
INIT_02 => X"918425005D45A411060604228642890040A491061E213031012C8000D7030206",
INIT_03 => X"6860699410016D322440A8D20600910304200004210010AA4082501400108001",
INIT_04 => X"AFFF9D8F603C2169A70150280207E432004880C5C0147145B1A0788B0638B911",
INIT_05 => X"C102609A62E44401230244A910230049482021090431009161FD24109000000A",
INIT_06 => X"C1BD40D46D080351A5B0A506EB684DD140BD0611E8998218802C8012C10401E9",
INIT_07 => X"A7056C8238820158E6980032BEB03FF08E21A02A2084008A18A3860404CD3890",
INIT_08 => X"2D89A40010321280520C894819004C070000C0B34342A4120901008001817B0A",
INIT_09 => X"0000000000000000005FFFFFFFFFFFEF7800000EF9FA8F76FC3ED7FDBCFDE954",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08C0708E06000000000000000D7FF80000FE01E94A845609155FFC000100002",
INIT_01 => X"081425AC41440812842012C018610038A10804B00C14A062001000C08000100C",
INIT_02 => X"120420020080A411054204280152000008809101410220044820000080210142",
INIT_03 => X"400010080000081208585489802024C014200004012E08805082000000121000",
INIT_04 => X"0000605096408404000A00000040142940480000000020810000104204100108",
INIT_05 => X"210A401822E44400980130A91038094040202CACA6804012000065CACAFA2240",
INIT_06 => X"040D0094000521402410040008082000481400034AE2420CA009801281040000",
INIT_07 => X"401004801002102384824420008081500401A48814A4200801010432B2801000",
INIT_08 => X"09802701C9F2130806EC804230180201000A03240039AA954AB4AA5085000B82",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE83BF7F7867CEE7F72EAD507FCFC7CF8A0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4CC031862648000000000000000000000000000840844008100000000100006",
INIT_01 => X"0804250020440802842102C012099610A10040B009001060000008C014000C2C",
INIT_02 => X"10040010008024110402040001D2040000809100410220144820000090210042",
INIT_03 => X"40001008001210084840108880600C4034200000000000098080000000100000",
INIT_04 => X"0000002080004802008608000140110048080000000228810004144205140428",
INIT_05 => X"4040401020E120828905102480A310501C10A02820C040020000000202000000",
INIT_06 => X"240D23F991019008240444040088200140148002A20082088008800000040026",
INIT_07 => X"00100481140A8081848A4220200884504503A06E068400280100800080009420",
INIT_08 => X"0264260101B1D102040428480810841500040002000030D86C382C1001000312",
INIT_09 => X"0000000000000000001FFFFFFFFFFFF200000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"D4C80010020C811111111111000000000000000000800C000100000000000002",
INIT_01 => X"0804258021440812842112C000099638A10844B000141062000009C814800C2C",
INIT_02 => X"100400100000A411040204200042000000801100400220140020000090010042",
INIT_03 => X"5000000808020A1000584481840028C204200004012E0888D080000000301000",
INIT_04 => X"A000621010418645C45946AAA800100900480002000004014000020204024000",
INIT_05 => X"210A400022240000190030A80019280048000C8C9210040280002DC84DFC22CA",
INIT_06 => X"00001050032460500004840000A8044040004009000002048008801281040024",
INIT_07 => X"0000048002000000848800202008001000810026506200040101963236C80210",
INIT_08 => X"141D0401CA5011080400000210180E010006400200191A0D068C864421000000",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE74B67630200DA6122CCA8C0FCFC7D6140",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100204811111111111000000000000000084084C008100000000100002",
INIT_01 => X"0010250AA0440812840112C000609228A10044B00000B060000008C014000C2C",
INIT_02 => X"B2042780008024110402040001D2046008C00001010264104A30200292214103",
INIT_03 => X"5000100808000A100850448800202C0014200004012E088050827814C2B20003",
INIT_04 => X"A000600010408441840142AAA840100900480002000102814002414204814008",
INIT_05 => X"A10A401822C440008001008900292840480024849280441280006D484DFC22CA",
INIT_06 => X"140908D0012420502404840400A825400004208848080204A0088012C1040000",
INIT_07 => X"021084808162102084880020200884502059842A50A420480100961212CA0110",
INIT_08 => X"0000260049E010000404804030080A00200A402200092A158A94CA4421000302",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE4234A4E04D5408102225FC4FD58D98220",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100264811111111111000000000000000084884C008100000000100002",
INIT_01 => X"0810250360440812840112C000609228A10044B00000B060000808C014000C2C",
INIT_02 => X"10040000000024110402040001520000008011010102201048200000D0210102",
INIT_03 => X"4000000800000810004800880020041014200000052C00805080000000100000",
INIT_04 => X"A000600010408441840142AAA800143000480000000100010002000204800000",
INIT_05 => X"C10A401222E40000810100A8003210484800280814C0400200002D8081BE224A",
INIT_06 => X"1489005002004010A0008404002025500804000808000208A0088052C1040000",
INIT_07 => X"4210008080020001048A4020200080402001800C00C400480101062024CA0010",
INIT_08 => X"0000260081B00080040401423010040100040002001030180C180C0001000302",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE771F0778E5016F81494EC15A01C5DA140",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C2880203B0600020202020200000000000400000000004001100000000000006",
INIT_01 => X"082425AC40448882840602C168004100A10180B0B4004064000000C00000000C",
INIT_02 => X"110400121014A411074204280042010000801104540220240024000080010042",
INIT_03 => X"40000888000041002040009302000181042000000000000A8080000000100000",
INIT_04 => X"0355134A4410692C60861400000010000008000080000B0100800582072A2001",
INIT_05 => X"0000400020000000320064000000000008000000000000022000000000000000",
INIT_06 => X"802050500000000100000400420000000029400000010200802D8000000400AC",
INIT_07 => X"8C0518832A800212449004200C200A20CA81008000000000010000000004AA00",
INIT_08 => X"0004050000000000040008080800801400000012002000000000000085030080",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE7394D4E04C1148010440605A158D94040",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C88A1F83F000020022002200020000000040004000000480012A000000000002",
INIT_01 => X"081025A00054C8C6940202C06F000801A50080B037810465AA0C60C00000008C",
INIT_02 => X"110400125014A4110746042880428100008411010603302100248000C0030106",
INIT_03 => X"4000018800010400044000DB822095C1142000002000102B8080000000100000",
INIT_04 => X"0F9B1B4E8208012E62940800020010000008808100000A4120000502072F8000",
INIT_05 => X"0040400260000001BA0374000000000808000000002100024000000000000000",
INIT_06 => X"81A078504000000180002502604008800029E01000000210802D8000000400EF",
INIT_07 => X"000400832F6000410692403298002000CBD90000000000A0012200000004AF80",
INIT_08 => X"0004070000001180040001000000000000000002400000000000000001806000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE701B2B18095005C029A93123518991024",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C6CC00100206811133331111580000000000010084084480A320000000100002",
INIT_01 => X"083425A020C40812840552811060DB28A10144A08801F060003809C014000C2C",
INIT_02 => X"114400321014A4110742042803520800408011054102201449240000D4210342",
INIT_03 => X"4800000800016D300048A0880020041014200001832C10A85080020000104400",
INIT_04 => X"ACE2ED56765C846DC75B56AAAA00109204480849C007540130A62A020480A800",
INIT_05 => X"410A401226C400218203048800321448480029091490400A60042D9091BE225A",
INIT_06 => X"7599005002184000A1002402434028800004001004000208800D8032810400E0",
INIT_07 => X"A515688080020959648240201830A2E02001820C20C4104A01030C2424820080",
INIT_08 => X"0004270091B0008034044140101044020004801A0052341A8D194C821101530A",
INIT_09 => X"0000000000000000005FFFFFFFFFFFF83800001EF9FE0F76FC3ED7DDE4E5F8C0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C088000001600222000000005A0000000040014000000480012A000000000002",
INIT_01 => X"08002500004408028400828000600000A10020A00000A060000000C00000000C",
INIT_02 => X"1084000000002411040204000042000000801100000220000028000081010002",
INIT_03 => X"4000000800000000004000800000000004200000000000000080000000108000",
INIT_04 => X"000D873106394000021014000200100000080000000000010000000204000000",
INIT_05 => X"0000400020000000000000000000000000000000000000020000000000000000",
INIT_06 => X"0000001000000000000004008000000000000000000002008008800000040000",
INIT_07 => X"0000008000000000048000200600000000010000000000000100000000000000",
INIT_08 => X"0000440000000000040000000000000000000002000000000000000001000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE07BF7F78E54CEFD36FAFD17FCFC7CF320",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08800000060022222222222000000000040000000000400010A000000000002",
INIT_01 => X"08002500004408028400028000000000A10000A000000060000800C00000000C",
INIT_02 => X"1004000000002411040204000042000000A01102160220000020000080010002",
INIT_03 => X"4000298800000000244008800000000004200000000000000080000000100000",
INIT_04 => X"0000008000042B24218800000200100000080000000001450000008A04000011",
INIT_05 => X"0000400020000000000000000000000000000000001000020000000000000000",
INIT_06 => X"0000001000000200002004000000000000000400000102008008800000040000",
INIT_07 => X"0000008000800000048000200000080000210000000000020100000000000000",
INIT_08 => X"0000040000001000040000000000000000000002000000000000000001000000",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"05104816EA00C199999999998B82D55555055577C0000675C3816AAAAAB80003",
INIT_01 => X"8014102000081213688B1862C400120ADA22C61962221218A90010E0957F0E0E",
INIT_02 => X"C200BAC50001061C8901300A2C0980A50085C801003641100400A00980206443",
INIT_03 => X"E2D5423CB284889002E20281C02900E8CC00000340A9401040162E6680824001",
INIT_04 => X"DAC651494D654F010FCA0208282AB2000D98181C14FDFC29876BFE33310017A2",
INIT_05 => X"0162E5846A0444221C5838881100401021048000000145D30AA9290000198B2F",
INIT_06 => X"84140A00A840000022800281241080040000104000002F219092A594094A9406",
INIT_07 => X"00000001010104011A42801D0244100440014000800490D0B58C444000A08004",
INIT_08 => X"612A8AB000AC00B4C66130400020000011002743150000000000100000548522",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE0334A4A0C60F6FB363875D4C538399B91",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4F74BF57E6E587FFFFFFFFFF92D71999998E665DC000E1D9E8758CCCCCF80000",
INIT_01 => X"2ADE30F033C915094A13393EDEF4B2265284CE4B6F40B85001AE0AB1FA003513",
INIT_02 => X"664123B786736A3991E3A47C1D59727F83855D59A1AC21CA6C30AAA2F8F149E3",
INIT_03 => X"01EF407061DE98DF4182021FC45117E22A0888D2C6F8E0FE6823B275CDE77725",
INIT_04 => X"D90A855E9396159B5AEBFD777C19EBC03DF139380EEDFC180363FE101FCE17A2",
INIT_05 => X"078D83F7F3CEFAFFFC5FFB96EBC021EE7D7ED00008BD6BB0067A7300009CCDED",
INIT_06 => X"5FEBF17BF430142FF1415AD12C11700001FFC007E7FAE8210DCA47FF1E58E6B8",
INIT_07 => X"105801B3FEE93C0112E1DACF82C6D945FFBB0E504085A1D076041DC000A6CE27",
INIT_08 => X"E66D1FC40024DFE9C023F3F007600088771815600D0020100800010630ECAF77",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE00C363180DDE2F82193AAC100343592A0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"80900040060040000000000040039E1E1E0F80060E1C067E2F81CF0F0F000003",
INIT_01 => X"82500F0000100211A6110064200002886984501A10005048A99041D0557F0A28",
INIT_02 => X"C0404B0000108804C04211220424A28000C0804940226454001080009001A502",
INIT_03 => X"6078001C3080000000EB02801129001CDC40000100810011D008380302004002",
INIT_04 => X"A662F955E7094500A5D54008A007F014021880C4040200098204001310000002",
INIT_05 => X"5062E0880ED505001C0038001036D20000002A1A1500108301F98CA1A12F1240",
INIT_06 => X"A4150A040AC0C8020A920A081014C00C2080386000000B2A5882A400218B3806",
INIT_07 => X"00500000008200051B06814AC10000000020810D82484020198561286D113146",
INIT_08 => X"266BAC10A190201046240000001405208005018303969048A41A4C084AD08000",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE00917109AA06CA940889D014484C5D990",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"00014020080007FFFFFFFFFF82D7E01FE008005FC000E7E1C1F5F00FF0380003",
INIT_01 => X"0000000000000004108800000000000104220004006A80000000000000000000",
INIT_02 => X"00009440000005400C0000020400000000000000002200000020000940000000",
INIT_03 => X"6040001C3080000000E20280000900000C000000000000000014440010000010",
INIT_04 => X"018F03201F7C056400DE0C82A800700000180004040000098200001310000002",
INIT_05 => X"0000E08000000000000000000000000000000000000000830018000000302240",
INIT_06 => X"000000000000000000000100000000000000000000000B20831BA40000240100",
INIT_07 => X"0000000000000000000000100000000000000000000000001184000000000000",
INIT_08 => X"2110402000000000462000000000000000000103010000000000000000000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE02EDADE84C87AAA0501480081CC8CB890",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"00000000000007FFFFFFFFFF82D7FFE0000FF85FC000E7E1C1F5FFF000380003",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000027C00000180004400007E00000000000000000000",
INIT_03 => X"E7C6867DF780000093E60380000900000C000000000000000000000000000000",
INIT_04 => X"A01182938901EA66400042A800BFF000001800043F10023B8E18013770310046",
INIT_05 => X"0000EF8000000000000000090000043020040000000007CF1FF800000401401A",
INIT_06 => X"000000000000000000000000000000000000000000001F200002A40000000000",
INIT_07 => X"00000004012900000000000000001004004B400000101001F99C000000000000",
INIT_08 => X"E0040100040C4805EEE00000000000000000230F3F0000000000112000000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE0402621121D803000120200200848E033",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4410801502168D555555555520D7FFFFFF90001F8000057F8D55FFFFFFF00002",
INIT_01 => X"8880BE000439376128C090A2E09240284A30242970600098540084F0017FA04B",
INIT_02 => X"0511481A600817F8800B64437D11428202208800047EF900C80488000085480F",
INIT_03 => X"E7D80EFFF7CC20E513E60BF2044D11000C800040108C0022022B789ECAA60068",
INIT_04 => X"A339708A60102128A000100000BFF000281B33343C01007B8E02003FFA280436",
INIT_05 => X"0400FF909010C50924424A0A4E0001004202001000202BC71FF8010000B8224A",
INIT_06 => X"803440026C000403008142D00504C00C20E91842A2A29FA1D882B4013A0BC088",
INIT_07 => X"21004806380200410AC4DA18814000418A00800040002047F9DC000040152848",
INIT_08 => X"F7F9E20001A3C285CFE02200024000A2D500B307BF0020100800000000F05610",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE038888C1EF9FE0FF6FC3CD7FDFCFD78DB",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"6CD0E84501520D555555555524FFFFFFFF90009F8001C17F8055FFFFFFF00000",
INIT_01 => X"0A94BEAFE77D3C314A43D337A45241685290F4CFD22090F85C488C03D57FAC62",
INIT_02 => X"F6157F9A78589FFDD14B756901537001E028C4415900AB14E83DA22A50A5694B",
INIT_03 => X"0827A802001090086000807A1124150890A222023DA002AA52AE78DFEAF6314B",
INIT_04 => X"AFBB390A30488569A60142AAAA0003022943B3B043B10100111A80008AA81AC0",
INIT_05 => X"052A101242D56D8BA4574A886E20405943422101103308000007AC10111C264A",
INIT_06 => X"95B9400000680303A0700FD92A012001036D0602A2A68081D98111502ADFFEA8",
INIT_07 => X"84170066A882B0892642407D02A2B185AA202C00A20445CC006054040096280A",
INIT_08 => X"17FD23001023D3900105A3409342604044500400800084422111088C6164DF12",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE07B77739EF5EEFB76BAFF15E4BCFDF3A8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"8A99D0720284A800000000006A000000005FFF400C1804002D00000000000002",
INIT_01 => X"A00080000420E3E7BC8241B640909201EF20906F206006E5F4E2B4F0200040CD",
INIT_02 => X"A39050087D451C8190084003FC04B16802C11910167EDC8180382AA20006800C",
INIT_03 => X"E7C02FFFF780000017EE0BA0044D00122CC888D0700CC010020D0094F2A38B73",
INIT_04 => X"0CCAAD86201C00280300100000BFF010001A02043C0C517F8E6028BFF0000017",
INIT_05 => X"4000FFC89801B282044400068092100014108808048043C71FFF818080920000",
INIT_06 => X"41040000420040000B034B10850100000010002000013FA88082B4013ADFFF40",
INIT_07 => X"000000000008000109A00A58044208000002004400420003FDFD002024201006",
INIT_08 => X"E000800080100005CFE00000001004A091043B97FF1200000008000002F83400",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE00000000000000000000000000000001B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010800820001080000840037C00000000000000007E88008380000000040008",
INIT_03 => X"E7C0067FF780000013E603A0000D00000C800000100000000210008001000040",
INIT_04 => X"0065E581003800000200100000BFF000001A02043C00003B8E000037F0000006",
INIT_05 => X"0000FF8000000000000000000000000000000000000003C71FFF800000300000",
INIT_06 => X"000000000000000000000000000000000000000000001FA00262B40281000000",
INIT_07 => X"000000000000000000000002400000000000000000000001F9DC000000000000",
INIT_08 => X"E000400000000005CFE000000000002091002307BF0000000000000000000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE01D1A18B4B598CC60523ACB39BEBD603B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010000820001080000840037C00028600040000007E88008000000000040008",
INIT_03 => X"E7D8067FF7DC38FD53E623A0000D00000C800000100000000200008000000040",
INIT_04 => X"0000600C600421202100000000BFF000001A02043C00203B8E001037F0100426",
INIT_05 => X"0000FF8000000000000000191120214040200010000027D71FFF890105B40080",
INIT_06 => X"0000032FBC009428008000005014C00C2080184000001FA00002B40000000000",
INIT_07 => X"A5414910100200586004900081100AE00400800840802001F9DC000040010060",
INIT_08 => X"E002201C05A0000DCFE00000002000229108A327BF0230180C100C0000002200",
INIT_09 => X"0000000000000000003FFFFFFFFFFFE020272920E9ED0B200C52CF20B83A81DB",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"85F820440E61E5DDDDDDDDDD81D7FFFFFF8FFE3FDEBCEF7FDFD5FFFFFFF80007",
INIT_01 => X"AA5E3FF033CC1A1BA4993AAC8064328EE9265EAA400ABA7000401AC1DE00573E",
INIT_02 => X"F645FFF78F73EF7DDDE3B57E7C6F72BF89C15D49E0FE675E24302AA9F8D1E5E3",
INIT_03 => X"E7FFD67DF7DE1ADFDBEF578C5479263E7E600053CEFDE25C78BFFE7FDFF77F3F",
INIT_04 => X"F000600019C294D19C21E3FFFDFFFBDD7FF9393C3FF980BB8F5BC0777CC057EE",
INIT_05 => X"76AFEFFFBFDFFFFEC44D899FFFFFFFFE7D7EFEBEBFDE7FFF1FFBFFEBEFFFFFFF",
INIT_06 => X"1ECB83FFBFF5FD6EFED75ED91C9CF11D68861AE7475A7F2FDFDBE7EFBFFFFF30",
INIT_07 => X"525A85B4C00BBCA59DE7DBED41CEC5553003EF7FD6FFF159FF9DFDFAFFB34067",
INIT_08 => X"FFFFFFFDEFFFFFFFEEEFF3F2377C0F29F31F676F3F9DBA9D6EAEBF7E7B7C8F77",
INIT_09 => X"0000000000000000003FFFFFFFFFFFE0034B422CD53444E373420BBD2C2CFAB3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"11200008002844CCCCCCCCCC80D7FFFFFF8FFE1F5AB4AB7F5ED5FFFFFFEA8015",
INIT_01 => X"080A0E5012800008002029000029049200080A4000142822000002090A800110",
INIT_02 => X"4441D8370DC3416110A004547C8854AB88011100A0FC000A040022202A1000A0",
INIT_03 => X"97EF9671EFDC1ADDDB97570404512A062A000057CA7F0844783D024B19456E38",
INIT_04 => X"F000600019C294D19C21E3FFFDFFEEED6471292A3FB880BA4F598074784056EE",
INIT_05 => X"B08F8FF597FFB2B2410480BECEADCE767554B6B6BBCC7BEC9FFBBF6B6BFDFF7F",
INIT_06 => X"0E4383AFBDD5BD7A76D7C05C1CACF55C688218EC0C023C267842452AEBF3DE10",
INIT_07 => X"5A189424400B2A2290A9DE0561CCC5511002CAEB96BD5119FE1CEE9ADBF94076",
INIT_08 => X"FFFF31FD6BEFE677E8EF78FA3E4C8B1D1113474C3F2DAA956AA6BB7AD42E0FD3",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE03F1110E441278421012A097022228883",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4128400000606088888888888000000000000000420526004380000000080003",
INIT_01 => X"220A20501184080808802A90006000C202200AA40000A820004A02822A004110",
INIT_02 => X"B24427A5000A440440A21114001A00002288C440A980220A0CA1088828B120A2",
INIT_03 => X"0000000000008000800100041110020C8222220186D182D428827A14E2B25403",
INIT_04 => X"50000000098210901820A155540009C40D2018180000A0000001100000500000",
INIT_05 => X"15A5002D0D0A4D38405082013104A72722261202091E1438000012202401D9B5",
INIT_06 => X"0A46800000B00800500004000001100103520206A6A480028100406810240010",
INIT_07 => X"104A014050019880140100200006500414006601401B30140200388809005000",
INIT_08 => X"0000D0E0240C34682002D2B0852621C8444918E8000400400012112631000041",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE02064636888C821822C1405C480005B40",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A5F0A0540E75C5DDDDDDDDDD81000000000FFE20C60C677EC3D5FFFFFFD80003",
INIT_01 => X"805E1FFFF1C81619E659392E8076B2AE79965E4B402AB858000A0A71FF7FBF3B",
INIT_02 => X"E240FFF78F72EB588DE1A03E016D627D81408809E0FE455E66100001F850C5E1",
INIT_03 => X"E037C67C104E00C793E9038C403806345E4000438F5D604C281FFE7FDFA35F3F",
INIT_04 => X"F0000000098210901820A15554BFFBD43EB9191C03F1A03B811BD0370CD013C6",
INIT_05 => X"5285E07FAFDEDDF4C409891B75D6B6EE3D3C5A0A0D9C1FFF0003F2A0A4BFFBFF",
INIT_06 => X"1ACE817992B0592EDA015AC90010100001160005455A5F0B5E9BE3FFAE2BE130",
INIT_07 => X"100800B0D0011C0519C74BCC4004400034014755405DB059FF813DE82D92502F",
INIT_08 => X"17FFDFE8A4BFFFEDEE03D1B0173405A8A20D37EF00941008040A15263A748175",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE0F480845EF1DE1EFDF8B9DEFDFCFDF890",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000222222222225A00000000000140000000800020000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE03B7F7BFCFDFCEFE37F7E0FFDBCBDF3E0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"60008010001404444444444400D7FFFFFF8FFE1F0810817F0C55FFFFFFE00000",
INIT_01 => X"08800E0FC20105004A40000200128020129000010020000800000030017FA801",
INIT_02 => X"4401D8120D410161100004407D1050EB80011110017C00804A00222200200800",
INIT_03 => X"87EF8671E7DC18DD5386030004410002280888D2492C0080503D004B19452A38",
INIT_04 => X"A000600010408441840142AAA8BFE200205121203FB8003A0F588034780016E6",
INIT_05 => X"010A8FD092D5B2820004009ECEA040505450A01010806BC41FFBAD0101BC264A",
INIT_06 => X"0401032FBC40952822D340581C04E00C20C0186000003C2058420512ABD3DE00",
INIT_07 => X"00100004000A200000A0DA0541C081410002884882844109F81C440040B1006C",
INIT_08 => X"F7FF211C01A3C215C8E5204012400000111007043F00A05028100808402C0F12",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE000000000000000000000000000000003",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA9918630DD2200000000000012800000040002000A106001180000000008003",
INIT_01 => X"80202100005CD2C7B4E6C1E566434955ED29B05AB311C477A91660C2B4D5208F",
INIT_02 => X"11840040D2AC24048604810082640D046B24CC461E01332121AD800087828206",
INIT_03 => X"080029800001E5202400B85242009129400A2A042000F22200808420C4108104",
INIT_04 => X"0FFF9D8F603C2128230010000300000242808041C004734430A038880239A811",
INIT_05 => X"020000002020000D274A4D200001018000080121202B00006004001212000000",
INIT_06 => X"C13448904109024705203C02E34808904139041A0823001024AC0285140000C9",
INIT_07 => X"AD0779C239A085FCE05801AA9E302EA48E692112240280820422814480043883",
INIT_08 => X"00008C001000080010000202A902E8120440D05040C204C2C131209008137028",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE0339694847C449F420A40C36848097824",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C084510228082000000000000020000000000000100004000108000000028006",
INIT_01 => X"22402100005000008490005046680400213C00142300E04080F4514BA066C00C",
INIT_02 => X"00000000000020044C00010000C28410230CC4480000024000A1800182C12400",
INIT_03 => X"00001000000000000810440001002000802880040000A2020000800004000000",
INIT_04 => X"006D858F60240028030010000140042911000040000032800000194004190008",
INIT_05 => X"A400000020200008014002200009080109000484820B00000000004848400000",
INIT_06 => X"010448504104201100008100002905400211220002A480048118000054040008",
INIT_07 => X"024205F019200280860000100002101406492022102200040000821212481910",
INIT_08 => X"080004204840000000080A08000A2A454002080000090A458294C24001820004",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE0614546024C1E10064251C088C4057AA0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0C0400000682101010101000092D555550554161001447421116AAAAA820012",
INIT_01 => X"0A001DAAA04408028418019800610454A10E00C4000CA262012000C8A0780028",
INIT_02 => X"100400120DC92A5D0C4335282951264102C1C140091444504A900282D2604003",
INIT_03 => X"82921220A28080400A92560001002012E062020401AE088010808000E4110B00",
INIT_04 => X"8000400010008001800040A2216AA439410080C0150120A80412106024900048",
INIT_05 => X"25280502622420C2000400A080C908191E12C4ACB24801600AA8284ACB6C0208",
INIT_06 => X"148401F4350564088D5442812C85210C221008A80880840DE318001020869400",
INIT_07 => X"025294C0908082810984424022C89D102421207614640008B4088012B2221060",
INIT_08 => X"4B3D0D0149D2C586804809008008A21544460200150B9A8D46B4AE500242A910",
INIT_09 => X"0000000000000000001FFFFFFFFFFFF62A53D68064DC5B30EAD404FCF071D0A1",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C081002008E009100110011024C366666619989C00210D460141B33333020006",
INIT_01 => X"0004B52CA4642830841112880080922C210C4480004812E055808C413181DC4C",
INIT_02 => X"101400182DD13AA94549640B18C2C44822849440480EA8148220888292050048",
INIT_03 => X"3183106A69989A5449B054A8102C240814A02200102C08101280808005100940",
INIT_04 => X"00000000104000410400408289599019410A02020D802098421090509410426A",
INIT_05 => X"E02873200000280081010000A00818001C0204ACA6C343038663254A4ACA200A",
INIT_06 => X"040C015D38052540005005141C14210422140822A0A429850A09B00002131800",
INIT_07 => X"0210048010000082068A043000C2811004010080142004006145001292801040",
INIT_08 => X"D19486014BD283038520180021088AD1514649018C298A8542BCAA5085880C80",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE450C1460054143016A2C000887031D238",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C48B20BC128580000111100000FC78787806181810000D18095E3C3C3C028006",
INIT_01 => X"0800252A604408128400100081842028A108042040C20260028008C0D0001E0C",
INIT_02 => X"920406120DD124110D42040879D2002022409100095E641048102008D2214003",
INIT_03 => X"87840669E7D0108253B6470800292C1018000000002E28001080601083130802",
INIT_04 => X"A00060000000000184010202A1B86529085010103E41203A0E02503474900026",
INIT_05 => X"60088F0A2A04610881110089810A09085C00048C828243571E19014848F0008A",
INIT_06 => X"1484017E820421508016840008A0A449401010C9832ADD24801B2400040C2100",
INIT_07 => X"0012848090001023048A4420008A9510240104A010202005E11C0612126A1010",
INIT_08 => X"DB9507014DC282878CE88108103AAE30F30E2B243C299A0D069C8E4085020880",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE949202102283E622408110054C4451803",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"CEC8381F030781111000000000D7807F8048181E94284D60B555C03FC0120006",
INIT_01 => X"082025836054C8D69416D281E46C6D2DA50DA4A0F217E665A82460C8448012AC",
INIT_02 => X"918425005D45A411060604228642890040A491061E213031012C8000D7030206",
INIT_03 => X"6860699410016D322440A8D20600910304200004210010AA4082501400108001",
INIT_04 => X"AFFF9D8F603C2169A70150280207E432004880C5C0147145B1A0788B0638B911",
INIT_05 => X"C102609A62E44401230244A910230049482021090431009161FD24109000000A",
INIT_06 => X"C1BD40D46D080351A5B0A506EB684DD140BD0611E8998218802C8012C10401E9",
INIT_07 => X"A7056C8238820158E6980032BEB03FF08E21A02A2084008A18A3860404CD3890",
INIT_08 => X"2D89A40010321280520C894819004C070000C0B34342A4120901008001817B0A",
INIT_09 => X"0000000000000000005FFFFFFFFFFFEF7800000EF9FA8F76FC3ED7FDBCFDE954",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08C0708E06000000000000000D7FF80000FE01E94A845609155FFC000100002",
INIT_01 => X"081425AC41440812842012C018610038A10804B00C14A062001000C08000100C",
INIT_02 => X"120420020080A411054204280152000008809101410220044820000080210142",
INIT_03 => X"400010080000081208585489802024C014200004012E08805082000000121000",
INIT_04 => X"0000605096408404000A00000040142940480000000020810000104204100108",
INIT_05 => X"210A401822E44400980130A91038094040202CACA6804012000065CACAFA2240",
INIT_06 => X"040D0094000521402410040008082000481400034AE2420CA009801281040000",
INIT_07 => X"401004801002102384824420008081500401A48814A4200801010432B2801000",
INIT_08 => X"09802701C9F2130806EC804230180201000A03240039AA954AB4AA5085000B82",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE83BF7F7867CEE7F72EAD507FCFC7CF8A0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4CC031862648000000000000000000000000000840844008100000000100006",
INIT_01 => X"0804250020440802842102C012099610A10040B009001060000008C014000C2C",
INIT_02 => X"10040010008024110402040001D2040000809100410220144820000090210042",
INIT_03 => X"40001008001210084840108880600C4034200000000000098080000000100000",
INIT_04 => X"0000002080004802008608000140110048080000000228810004144205140428",
INIT_05 => X"4040401020E120828905102480A310501C10A02820C040020000000202000000",
INIT_06 => X"240D23F991019008240444040088200140148002A20082088008800000040026",
INIT_07 => X"00100481140A8081848A4220200884504503A06E068400280100800080009420",
INIT_08 => X"0264260101B1D102040428480810841500040002000030D86C382C1001000312",
INIT_09 => X"0000000000000000001FFFFFFFFFFFF200000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"D4C80010020C811111111111000000000000000000800C000100000000000002",
INIT_01 => X"0804258021440812842112C000099638A10844B000141062000009C814800C2C",
INIT_02 => X"100400100000A411040204200042000000801100400220140020000090010042",
INIT_03 => X"5000000808020A1000584481840028C204200004012E0888D080000000301000",
INIT_04 => X"A000621010418645C45946AAA800100900480002000004014000020204024000",
INIT_05 => X"210A400022240000190030A80019280048000C8C9210040280002DC84DFC22CA",
INIT_06 => X"00001050032460500004840000A8044040004009000002048008801281040024",
INIT_07 => X"0000048002000000848800202008001000810026506200040101963236C80210",
INIT_08 => X"141D0401CA5011080400000210180E010006400200191A0D068C864421000000",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE74B67630200DA6122CCA8C0FCFC7D6140",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100204811111111111000000000000000084084C008100000000100002",
INIT_01 => X"0010250AA0440812840112C000609228A10044B00000B060000008C014000C2C",
INIT_02 => X"B2042780008024110402040001D2046008C00001010264104A30200292214103",
INIT_03 => X"5000100808000A100850448800202C0014200004012E088050827814C2B20003",
INIT_04 => X"A000600010408441840142AAA840100900480002000102814002414204814008",
INIT_05 => X"A10A401822C440008001008900292840480024849280441280006D484DFC22CA",
INIT_06 => X"140908D0012420502404840400A825400004208848080204A0088012C1040000",
INIT_07 => X"021084808162102084880020200884502059842A50A420480100961212CA0110",
INIT_08 => X"0000260049E010000404804030080A00200A402200092A158A94CA4421000302",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE4234A4E04D5408102225FC4FD58D98220",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100264811111111111000000000000000084884C008100000000100002",
INIT_01 => X"0810250360440812840112C000609228A10044B00000B060000808C014000C2C",
INIT_02 => X"10040000000024110402040001520000008011010102201048200000D0210102",
INIT_03 => X"4000000800000810004800880020041014200000052C00805080000000100000",
INIT_04 => X"A000600010408441840142AAA800143000480000000100010002000204800000",
INIT_05 => X"C10A401222E40000810100A8003210484800280814C0400200002D8081BE224A",
INIT_06 => X"1489005002004010A0008404002025500804000808000208A0088052C1040000",
INIT_07 => X"4210008080020001048A4020200080402001800C00C400480101062024CA0010",
INIT_08 => X"0000260081B00080040401423010040100040002001030180C180C0001000302",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE771F0778E5016F81494EC15A01C5DA140",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C2880203B0600020202020200000000000400000000004001100000000000006",
INIT_01 => X"082425AC40448882840602C168004100A10180B0B4004064000000C00000000C",
INIT_02 => X"110400121014A411074204280042010000801104540220240024000080010042",
INIT_03 => X"40000888000041002040009302000181042000000000000A8080000000100000",
INIT_04 => X"0355134A4410692C60861400000010000008000080000B0100800582072A2001",
INIT_05 => X"0000400020000000320064000000000008000000000000022000000000000000",
INIT_06 => X"802050500000000100000400420000000029400000010200802D8000000400AC",
INIT_07 => X"8C0518832A800212449004200C200A20CA81008000000000010000000004AA00",
INIT_08 => X"0004050000000000040008080800801400000012002000000000000085030080",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE7394D4E04C1148010440605A158D94040",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C88A1F83F000020022002200020000000040004000000480012A000000000002",
INIT_01 => X"081025A00054C8C6940202C06F000801A50080B037810465AA0C60C00000008C",
INIT_02 => X"110400125014A4110746042880428100008411010603302100248000C0030106",
INIT_03 => X"4000018800010400044000DB822095C1142000002000102B8080000000100000",
INIT_04 => X"0F9B1B4E8208012E62940800020010000008808100000A4120000502072F8000",
INIT_05 => X"0040400260000001BA0374000000000808000000002100024000000000000000",
INIT_06 => X"81A078504000000180002502604008800029E01000000210802D8000000400EF",
INIT_07 => X"000400832F6000410692403298002000CBD90000000000A0012200000004AF80",
INIT_08 => X"0004070000001180040001000000000000000002400000000000000001806000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE701B2B18095005C029A93123518991024",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C6CC00100206811133331111580000000000010084084480A320000000100002",
INIT_01 => X"083425A020C40812840552811060DB28A10144A08801F060003809C014000C2C",
INIT_02 => X"114400321014A4110742042803520800408011054102201449240000D4210342",
INIT_03 => X"4800000800016D300048A0880020041014200001832C10A85080020000104400",
INIT_04 => X"ACE2ED56765C846DC75B56AAAA00109204480849C007540130A62A020480A800",
INIT_05 => X"410A401226C400218203048800321448480029091490400A60042D9091BE225A",
INIT_06 => X"7599005002184000A1002402434028800004001004000208800D8032810400E0",
INIT_07 => X"A515688080020959648240201830A2E02001820C20C4104A01030C2424820080",
INIT_08 => X"0004270091B0008034044140101044020004801A0052341A8D194C821101530A",
INIT_09 => X"0000000000000000005FFFFFFFFFFFF83800001EF9FE0F76FC3ED7DDE4E5F8C0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C088000001600222000000005A0000000040014000000480012A000000000002",
INIT_01 => X"08002500004408028400828000600000A10020A00000A060000000C00000000C",
INIT_02 => X"1084000000002411040204000042000000801100000220000028000081010002",
INIT_03 => X"4000000800000000004000800000000004200000000000000080000000108000",
INIT_04 => X"000D873106394000021014000200100000080000000000010000000204000000",
INIT_05 => X"0000400020000000000000000000000000000000000000020000000000000000",
INIT_06 => X"0000001000000000000004008000000000000000000002008008800000040000",
INIT_07 => X"0000008000000000048000200600000000010000000000000100000000000000",
INIT_08 => X"0000440000000000040000000000000000000002000000000000000001000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE07BF7F78E54CEFD36FAFD17FCFC7CF320",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08800000060022222222222000000000040000000000400010A000000000002",
INIT_01 => X"08002500004408028400028000000000A10000A000000060000800C00000000C",
INIT_02 => X"1004000000002411040204000042000000A01102160220000020000080010002",
INIT_03 => X"4000298800000000244008800000000004200000000000000080000000100000",
INIT_04 => X"0000008000042B24218800000200100000080000000001450000008A04000011",
INIT_05 => X"0000400020000000000000000000000000000000001000020000000000000000",
INIT_06 => X"0000001000000200002004000000000000000400000102008008800000040000",
INIT_07 => X"0000008000800000048000200000080000210000000000020100000000000000",
INIT_08 => X"0000040000001000040000000000000000000002000000000000000001000000",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"05104816EA00C199999999998B82D55555055577C0000675C3816AAAAAB80003",
INIT_01 => X"8014102000081213688B1862C400120ADA22C61962221218A90010E0957F0E0E",
INIT_02 => X"C200BAC50001061C8901300A2C0980A50085C801003641100400A00980206443",
INIT_03 => X"E2D5423CB284889002E20281C02900E8CC00000340A9401040162E6680824001",
INIT_04 => X"DAC651494D654F010FCA0208282AB2000D98181C14FDFC29876BFE33310017A2",
INIT_05 => X"0162E5846A0444221C5838881100401021048000000145D30AA9290000198B2F",
INIT_06 => X"84140A00A840000022800281241080040000104000002F219092A594094A9406",
INIT_07 => X"00000001010104011A42801D0244100440014000800490D0B58C444000A08004",
INIT_08 => X"612A8AB000AC00B4C66130400020000011002743150000000000100000548522",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE0334A4A0C60F6FB363875D4C538399B91",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4F74BF57E6E587FFFFFFFFFF92D71999998E665DC000E1D9E8758CCCCCF80000",
INIT_01 => X"2ADE30F033C915094A13393EDEF4B2265284CE4B6F40B85001AE0AB1FA003513",
INIT_02 => X"664123B786736A3991E3A47C1D59727F83855D59A1AC21CA6C30AAA2F8F149E3",
INIT_03 => X"01EF407061DE98DF4182021FC45117E22A0888D2C6F8E0FE6823B275CDE77725",
INIT_04 => X"D90A855E9396159B5AEBFD777C19EBC03DF139380EEDFC180363FE101FCE17A2",
INIT_05 => X"078D83F7F3CEFAFFFC5FFB96EBC021EE7D7ED00008BD6BB0067A7300009CCDED",
INIT_06 => X"5FEBF17BF430142FF1415AD12C11700001FFC007E7FAE8210DCA47FF1E58E6B8",
INIT_07 => X"105801B3FEE93C0112E1DACF82C6D945FFBB0E504085A1D076041DC000A6CE27",
INIT_08 => X"E66D1FC40024DFE9C023F3F007600088771815600D0020100800010630ECAF77",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE00C363180DDE2F82193AAC100343592A0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"80900040060040000000000040039E1E1E0F80060E1C067E2F81CF0F0F000003",
INIT_01 => X"82500F0000100211A6110064200002886984501A10005048A99041D0557F0A28",
INIT_02 => X"C0404B0000108804C04211220424A28000C0804940226454001080009001A502",
INIT_03 => X"6078001C3080000000EB02801129001CDC40000100810011D008380302004002",
INIT_04 => X"A662F955E7094500A5D54008A007F014021880C4040200098204001310000002",
INIT_05 => X"5062E0880ED505001C0038001036D20000002A1A1500108301F98CA1A12F1240",
INIT_06 => X"A4150A040AC0C8020A920A081014C00C2080386000000B2A5882A400218B3806",
INIT_07 => X"00500000008200051B06814AC10000000020810D82484020198561286D113146",
INIT_08 => X"266BAC10A190201046240000001405208005018303969048A41A4C084AD08000",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE00917109AA06CA940889D014484C5D990",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"00014020080007FFFFFFFFFF82D7E01FE008005FC000E7E1C1F5F00FF0380003",
INIT_01 => X"0000000000000004108800000000000104220004006A80000000000000000000",
INIT_02 => X"00009440000005400C0000020400000000000000002200000020000940000000",
INIT_03 => X"6040001C3080000000E20280000900000C000000000000000014440010000010",
INIT_04 => X"018F03201F7C056400DE0C82A800700000180004040000098200001310000002",
INIT_05 => X"0000E08000000000000000000000000000000000000000830018000000302240",
INIT_06 => X"000000000000000000000100000000000000000000000B20831BA40000240100",
INIT_07 => X"0000000000000000000000100000000000000000000000001184000000000000",
INIT_08 => X"2110402000000000462000000000000000000103010000000000000000000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE02EDADE84C87AAA0501480081CC8CB890",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"00000000000007FFFFFFFFFF82D7FFE0000FF85FC000E7E1C1F5FFF000380003",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000027C00000180004400007E00000000000000000000",
INIT_03 => X"E7C6867DF780000093E60380000900000C000000000000000000000000000000",
INIT_04 => X"A01182938901EA66400042A800BFF000001800043F10023B8E18013770310046",
INIT_05 => X"0000EF8000000000000000090000043020040000000007CF1FF800000401401A",
INIT_06 => X"000000000000000000000000000000000000000000001F200002A40000000000",
INIT_07 => X"00000004012900000000000000001004004B400000101001F99C000000000000",
INIT_08 => X"E0040100040C4805EEE00000000000000000230F3F0000000000112000000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE0402621121D803000120200200848E033",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4410801502168D555555555520D7FFFFFF90001F8000057F8D55FFFFFFF00002",
INIT_01 => X"8880BE000439376128C090A2E09240284A30242970600098540084F0017FA04B",
INIT_02 => X"0511481A600817F8800B64437D11428202208800047EF900C80488000085480F",
INIT_03 => X"E7D80EFFF7CC20E513E60BF2044D11000C800040108C0022022B789ECAA60068",
INIT_04 => X"A339708A60102128A000100000BFF000281B33343C01007B8E02003FFA280436",
INIT_05 => X"0400FF909010C50924424A0A4E0001004202001000202BC71FF8010000B8224A",
INIT_06 => X"803440026C000403008142D00504C00C20E91842A2A29FA1D882B4013A0BC088",
INIT_07 => X"21004806380200410AC4DA18814000418A00800040002047F9DC000040152848",
INIT_08 => X"F7F9E20001A3C285CFE02200024000A2D500B307BF0020100800000000F05610",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE038888C1EF9FE0FF6FC3CD7FDFCFD78DB",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"6CD0E84501520D555555555524FFFFFFFF90009F8001C17F8055FFFFFFF00000",
INIT_01 => X"0A94BEAFE77D3C314A43D337A45241685290F4CFD22090F85C488C03D57FAC62",
INIT_02 => X"F6157F9A78589FFDD14B756901537001E028C4415900AB14E83DA22A50A5694B",
INIT_03 => X"0827A802001090086000807A1124150890A222023DA002AA52AE78DFEAF6314B",
INIT_04 => X"AFBB390A30488569A60142AAAA0003022943B3B043B10100111A80008AA81AC0",
INIT_05 => X"052A101242D56D8BA4574A886E20405943422101103308000007AC10111C264A",
INIT_06 => X"95B9400000680303A0700FD92A012001036D0602A2A68081D98111502ADFFEA8",
INIT_07 => X"84170066A882B0892642407D02A2B185AA202C00A20445CC006054040096280A",
INIT_08 => X"17FD23001023D3900105A3409342604044500400800084422111088C6164DF12",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE07B77739EF5EEFB76BAFF15E4BCFDF3A8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"8A99D0720284A800000000006A000000005FFF400C1804002D00000000000002",
INIT_01 => X"A00080000420E3E7BC8241B640909201EF20906F206006E5F4E2B4F0200040CD",
INIT_02 => X"A39050087D451C8190084003FC04B16802C11910167EDC8180382AA20006800C",
INIT_03 => X"E7C02FFFF780000017EE0BA0044D00122CC888D0700CC010020D0094F2A38B73",
INIT_04 => X"0CCAAD86201C00280300100000BFF010001A02043C0C517F8E6028BFF0000017",
INIT_05 => X"4000FFC89801B282044400068092100014108808048043C71FFF818080920000",
INIT_06 => X"41040000420040000B034B10850100000010002000013FA88082B4013ADFFF40",
INIT_07 => X"000000000008000109A00A58044208000002004400420003FDFD002024201006",
INIT_08 => X"E000800080100005CFE00000001004A091043B97FF1200000008000002F83400",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE00000000000000000000000000000001B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010800820001080000840037C00000000000000007E88008380000000040008",
INIT_03 => X"E7C0067FF780000013E603A0000D00000C800000100000000210008001000040",
INIT_04 => X"0065E581003800000200100000BFF000001A02043C00003B8E000037F0000006",
INIT_05 => X"0000FF8000000000000000000000000000000000000003C71FFF800000300000",
INIT_06 => X"000000000000000000000000000000000000000000001FA00262B40281000000",
INIT_07 => X"000000000000000000000002400000000000000000000001F9DC000000000000",
INIT_08 => X"E000400000000005CFE000000000002091002307BF0000000000000000000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE01D1A18B4B598CC60523ACB39BEBD603B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010000820001080000840037C00028600040000007E88008000000000040008",
INIT_03 => X"E7D8067FF7DC38FD53E623A0000D00000C800000100000000200008000000040",
INIT_04 => X"0000600C600421202100000000BFF000001A02043C00203B8E001037F0100426",
INIT_05 => X"0000FF8000000000000000191120214040200010000027D71FFF890105B40080",
INIT_06 => X"0000032FBC009428008000005014C00C2080184000001FA00002B40000000000",
INIT_07 => X"A5414910100200586004900081100AE00400800840802001F9DC000040010060",
INIT_08 => X"E002201C05A0000DCFE00000002000229108A327BF0230180C100C0000002200",
INIT_09 => X"0000000000000000003FFFFFFFFFFFE020272920E9ED0B200C52CF20B83A81DB",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"85F820440E61E5DDDDDDDDDD81D7FFFFFF8FFE3FDEBCEF7FDFD5FFFFFFF80007",
INIT_01 => X"AA5E3FF033CC1A1BA4993AAC8064328EE9265EAA400ABA7000401AC1DE00573E",
INIT_02 => X"F645FFF78F73EF7DDDE3B57E7C6F72BF89C15D49E0FE675E24302AA9F8D1E5E3",
INIT_03 => X"E7FFD67DF7DE1ADFDBEF578C5479263E7E600053CEFDE25C78BFFE7FDFF77F3F",
INIT_04 => X"F000600019C294D19C21E3FFFDFFFBDD7FF9393C3FF980BB8F5BC0777CC057EE",
INIT_05 => X"76AFEFFFBFDFFFFEC44D899FFFFFFFFE7D7EFEBEBFDE7FFF1FFBFFEBEFFFFFFF",
INIT_06 => X"1ECB83FFBFF5FD6EFED75ED91C9CF11D68861AE7475A7F2FDFDBE7EFBFFFFF30",
INIT_07 => X"525A85B4C00BBCA59DE7DBED41CEC5553003EF7FD6FFF159FF9DFDFAFFB34067",
INIT_08 => X"FFFFFFFDEFFFFFFFEEEFF3F2377C0F29F31F676F3F9DBA9D6EAEBF7E7B7C8F77",
INIT_09 => X"0000000000000000003FFFFFFFFFFFE0034B422CD53444E373420BBD2C2CFAB3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"11200008002844CCCCCCCCCC80D7FFFFFF8FFE1F5AB4AB7F5ED5FFFFFFEA8015",
INIT_01 => X"080A0E5012800008002029000029049200080A4000142822000002090A800110",
INIT_02 => X"4441D8370DC3416110A004547C8854AB88011100A0FC000A040022202A1000A0",
INIT_03 => X"97EF9671EFDC1ADDDB97570404512A062A000057CA7F0844783D024B19456E38",
INIT_04 => X"F000600019C294D19C21E3FFFDFFEEED6471292A3FB880BA4F598074784056EE",
INIT_05 => X"B08F8FF597FFB2B2410480BECEADCE767554B6B6BBCC7BEC9FFBBF6B6BFDFF7F",
INIT_06 => X"0E4383AFBDD5BD7A76D7C05C1CACF55C688218EC0C023C267842452AEBF3DE10",
INIT_07 => X"5A189424400B2A2290A9DE0561CCC5511002CAEB96BD5119FE1CEE9ADBF94076",
INIT_08 => X"FFFF31FD6BEFE677E8EF78FA3E4C8B1D1113474C3F2DAA956AA6BB7AD42E0FD3",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE03F1110E441278421012A097022228883",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4128400000606088888888888000000000000000420526004380000000080003",
INIT_01 => X"220A20501184080808802A90006000C202200AA40000A820004A02822A004110",
INIT_02 => X"B24427A5000A440440A21114001A00002288C440A980220A0CA1088828B120A2",
INIT_03 => X"0000000000008000800100041110020C8222220186D182D428827A14E2B25403",
INIT_04 => X"50000000098210901820A155540009C40D2018180000A0000001100000500000",
INIT_05 => X"15A5002D0D0A4D38405082013104A72722261202091E1438000012202401D9B5",
INIT_06 => X"0A46800000B00800500004000001100103520206A6A480028100406810240010",
INIT_07 => X"104A014050019880140100200006500414006601401B30140200388809005000",
INIT_08 => X"0000D0E0240C34682002D2B0852621C8444918E8000400400012112631000041",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE02064636888C821822C1405C480005B40",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A5F0A0540E75C5DDDDDDDDDD81000000000FFE20C60C677EC3D5FFFFFFD80003",
INIT_01 => X"805E1FFFF1C81619E659392E8076B2AE79965E4B402AB858000A0A71FF7FBF3B",
INIT_02 => X"E240FFF78F72EB588DE1A03E016D627D81408809E0FE455E66100001F850C5E1",
INIT_03 => X"E037C67C104E00C793E9038C403806345E4000438F5D604C281FFE7FDFA35F3F",
INIT_04 => X"F0000000098210901820A15554BFFBD43EB9191C03F1A03B811BD0370CD013C6",
INIT_05 => X"5285E07FAFDEDDF4C409891B75D6B6EE3D3C5A0A0D9C1FFF0003F2A0A4BFFBFF",
INIT_06 => X"1ACE817992B0592EDA015AC90010100001160005455A5F0B5E9BE3FFAE2BE130",
INIT_07 => X"100800B0D0011C0519C74BCC4004400034014755405DB059FF813DE82D92502F",
INIT_08 => X"17FFDFE8A4BFFFEDEE03D1B0173405A8A20D37EF00941008040A15263A748175",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE0F480845EF1DE1EFDF8B9DEFDFCFDF890",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000222222222225A00000000000140000000800020000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE03B7F7BFCFDFCEFE37F7E0FFDBCBDF3E0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"60008010001404444444444400D7FFFFFF8FFE1F0810817F0C55FFFFFFE00000",
INIT_01 => X"08800E0FC20105004A40000200128020129000010020000800000030017FA801",
INIT_02 => X"4401D8120D410161100004407D1050EB80011110017C00804A00222200200800",
INIT_03 => X"87EF8671E7DC18DD5386030004410002280888D2492C0080503D004B19452A38",
INIT_04 => X"A000600010408441840142AAA8BFE200205121203FB8003A0F588034780016E6",
INIT_05 => X"010A8FD092D5B2820004009ECEA040505450A01010806BC41FFBAD0101BC264A",
INIT_06 => X"0401032FBC40952822D340581C04E00C20C0186000003C2058420512ABD3DE00",
INIT_07 => X"00100004000A200000A0DA0541C081410002884882844109F81C440040B1006C",
INIT_08 => X"F7FF211C01A3C215C8E5204012400000111007043F00A05028100808402C0F12",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE000000000000000000000000000000003",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA9918630DD2200000000000012800000040002000A106001180000000008003",
INIT_01 => X"80202100005CD2C7B4E6C1E566434955ED29B05AB311C477A91660C2B4D5208F",
INIT_02 => X"11840040D2AC24048604810082640D046B24CC461E01332121AD800087828206",
INIT_03 => X"080029800001E5202400B85242009129400A2A042000F22200808420C4108104",
INIT_04 => X"0FFF9D8F603C2128230010000300000242808041C004734430A038880239A811",
INIT_05 => X"020000002020000D274A4D200001018000080121202B00006004001212000000",
INIT_06 => X"C13448904109024705203C02E34808904139041A0823001024AC0285140000C9",
INIT_07 => X"AD0779C239A085FCE05801AA9E302EA48E692112240280820422814480043883",
INIT_08 => X"00008C001000080010000202A902E8120440D05040C204C2C131209008137028",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE0339694847C449F420A40C36848097824",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C084510228082000000000000020000000000000100004000108000000028006",
INIT_01 => X"22402100005000008490005046680400213C00142300E04080F4514BA066C00C",
INIT_02 => X"00000000000020044C00010000C28410230CC4480000024000A1800182C12400",
INIT_03 => X"00001000000000000810440001002000802880040000A2020000800004000000",
INIT_04 => X"006D858F60240028030010000140042911000040000032800000194004190008",
INIT_05 => X"A400000020200008014002200009080109000484820B00000000004848400000",
INIT_06 => X"010448504104201100008100002905400211220002A480048118000054040008",
INIT_07 => X"024205F019200280860000100002101406492022102200040000821212481910",
INIT_08 => X"080004204840000000080A08000A2A454002080000090A458294C24001820004",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE0614546024C1E10064251C088C4057AA0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0C0400000682101010101000092D555550554161001447421116AAAAA820012",
INIT_01 => X"0A001DAAA04408028418019800610454A10E00C4000CA262012000C8A0780028",
INIT_02 => X"100400120DC92A5D0C4335282951264102C1C140091444504A900282D2604003",
INIT_03 => X"82921220A28080400A92560001002012E062020401AE088010808000E4110B00",
INIT_04 => X"8000400010008001800040A2216AA439410080C0150120A80412106024900048",
INIT_05 => X"25280502622420C2000400A080C908191E12C4ACB24801600AA8284ACB6C0208",
INIT_06 => X"148401F4350564088D5442812C85210C221008A80880840DE318001020869400",
INIT_07 => X"025294C0908082810984424022C89D102421207614640008B4088012B2221060",
INIT_08 => X"4B3D0D0149D2C586804809008008A21544460200150B9A8D46B4AE500242A910",
INIT_09 => X"0000000000000000001FFFFFFFFFFFF62A53D68064DC5B30EAD404FCF071D0A1",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C081002008E009100110011024C366666619989C00210D460141B33333020006",
INIT_01 => X"0004B52CA4642830841112880080922C210C4480004812E055808C413181DC4C",
INIT_02 => X"101400182DD13AA94549640B18C2C44822849440480EA8148220888292050048",
INIT_03 => X"3183106A69989A5449B054A8102C240814A02200102C08101280808005100940",
INIT_04 => X"00000000104000410400408289599019410A02020D802098421090509410426A",
INIT_05 => X"E02873200000280081010000A00818001C0204ACA6C343038663254A4ACA200A",
INIT_06 => X"040C015D38052540005005141C14210422140822A0A429850A09B00002131800",
INIT_07 => X"0210048010000082068A043000C2811004010080142004006145001292801040",
INIT_08 => X"D19486014BD283038520180021088AD1514649018C298A8542BCAA5085880C80",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE450C1460054143016A2C000887031D238",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C48B20BC128580000111100000FC78787806181810000D18095E3C3C3C028006",
INIT_01 => X"0800252A604408128400100081842028A108042040C20260028008C0D0001E0C",
INIT_02 => X"920406120DD124110D42040879D2002022409100095E641048102008D2214003",
INIT_03 => X"87840669E7D0108253B6470800292C1018000000002E28001080601083130802",
INIT_04 => X"A00060000000000184010202A1B86529085010103E41203A0E02503474900026",
INIT_05 => X"60088F0A2A04610881110089810A09085C00048C828243571E19014848F0008A",
INIT_06 => X"1484017E820421508016840008A0A449401010C9832ADD24801B2400040C2100",
INIT_07 => X"0012848090001023048A4420008A9510240104A010202005E11C0612126A1010",
INIT_08 => X"DB9507014DC282878CE88108103AAE30F30E2B243C299A0D069C8E4085020880",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE949202102283E622408110054C4451803",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"CEC8381F030781111000000000D7807F8048181E94284D60B555C03FC0120006",
INIT_01 => X"082025836054C8D69416D281E46C6D2DA50DA4A0F217E665A82460C8448012AC",
INIT_02 => X"918425005D45A411060604228642890040A491061E213031012C8000D7030206",
INIT_03 => X"6860699410016D322440A8D20600910304200004210010AA4082501400108001",
INIT_04 => X"AFFF9D8F603C2169A70150280207E432004880C5C0147145B1A0788B0638B911",
INIT_05 => X"C102609A62E44401230244A910230049482021090431009161FD24109000000A",
INIT_06 => X"C1BD40D46D080351A5B0A506EB684DD140BD0611E8998218802C8012C10401E9",
INIT_07 => X"A7056C8238820158E6980032BEB03FF08E21A02A2084008A18A3860404CD3890",
INIT_08 => X"2D89A40010321280520C894819004C070000C0B34342A4120901008001817B0A",
INIT_09 => X"0000000000000000005FFFFFFFFFFFEF7800000EF9FA8F76FC3ED7FDBCFDE954",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08C0708E06000000000000000D7FF80000FE01E94A845609155FFC000100002",
INIT_01 => X"081425AC41440812842012C018610038A10804B00C14A062001000C08000100C",
INIT_02 => X"120420020080A411054204280152000008809101410220044820000080210142",
INIT_03 => X"400010080000081208585489802024C014200004012E08805082000000121000",
INIT_04 => X"0000605096408404000A00000040142940480000000020810000104204100108",
INIT_05 => X"210A401822E44400980130A91038094040202CACA6804012000065CACAFA2240",
INIT_06 => X"040D0094000521402410040008082000481400034AE2420CA009801281040000",
INIT_07 => X"401004801002102384824420008081500401A48814A4200801010432B2801000",
INIT_08 => X"09802701C9F2130806EC804230180201000A03240039AA954AB4AA5085000B82",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE83BF7F7867CEE7F72EAD507FCFC7CF8A0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4CC031862648000000000000000000000000000840844008100000000100006",
INIT_01 => X"0804250020440802842102C012099610A10040B009001060000008C014000C2C",
INIT_02 => X"10040010008024110402040001D2040000809100410220144820000090210042",
INIT_03 => X"40001008001210084840108880600C4034200000000000098080000000100000",
INIT_04 => X"0000002080004802008608000140110048080000000228810004144205140428",
INIT_05 => X"4040401020E120828905102480A310501C10A02820C040020000000202000000",
INIT_06 => X"240D23F991019008240444040088200140148002A20082088008800000040026",
INIT_07 => X"00100481140A8081848A4220200884504503A06E068400280100800080009420",
INIT_08 => X"0264260101B1D102040428480810841500040002000030D86C382C1001000312",
INIT_09 => X"0000000000000000001FFFFFFFFFFFF200000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"D4C80010020C811111111111000000000000000000800C000100000000000002",
INIT_01 => X"0804258021440812842112C000099638A10844B000141062000009C814800C2C",
INIT_02 => X"100400100000A411040204200042000000801100400220140020000090010042",
INIT_03 => X"5000000808020A1000584481840028C204200004012E0888D080000000301000",
INIT_04 => X"A000621010418645C45946AAA800100900480002000004014000020204024000",
INIT_05 => X"210A400022240000190030A80019280048000C8C9210040280002DC84DFC22CA",
INIT_06 => X"00001050032460500004840000A8044040004009000002048008801281040024",
INIT_07 => X"0000048002000000848800202008001000810026506200040101963236C80210",
INIT_08 => X"141D0401CA5011080400000210180E010006400200191A0D068C864421000000",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE74B67630200DA6122CCA8C0FCFC7D6140",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100204811111111111000000000000000084084C008100000000100002",
INIT_01 => X"0010250AA0440812840112C000609228A10044B00000B060000008C014000C2C",
INIT_02 => X"B2042780008024110402040001D2046008C00001010264104A30200292214103",
INIT_03 => X"5000100808000A100850448800202C0014200004012E088050827814C2B20003",
INIT_04 => X"A000600010408441840142AAA840100900480002000102814002414204814008",
INIT_05 => X"A10A401822C440008001008900292840480024849280441280006D484DFC22CA",
INIT_06 => X"140908D0012420502404840400A825400004208848080204A0088012C1040000",
INIT_07 => X"021084808162102084880020200884502059842A50A420480100961212CA0110",
INIT_08 => X"0000260049E010000404804030080A00200A402200092A158A94CA4421000302",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE4234A4E04D5408102225FC4FD58D98220",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100264811111111111000000000000000084884C008100000000100002",
INIT_01 => X"0810250360440812840112C000609228A10044B00000B060000808C014000C2C",
INIT_02 => X"10040000000024110402040001520000008011010102201048200000D0210102",
INIT_03 => X"4000000800000810004800880020041014200000052C00805080000000100000",
INIT_04 => X"A000600010408441840142AAA800143000480000000100010002000204800000",
INIT_05 => X"C10A401222E40000810100A8003210484800280814C0400200002D8081BE224A",
INIT_06 => X"1489005002004010A0008404002025500804000808000208A0088052C1040000",
INIT_07 => X"4210008080020001048A4020200080402001800C00C400480101062024CA0010",
INIT_08 => X"0000260081B00080040401423010040100040002001030180C180C0001000302",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE771F0778E5016F81494EC15A01C5DA140",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C2880203B0600020202020200000000000400000000004001100000000000006",
INIT_01 => X"082425AC40448882840602C168004100A10180B0B4004064000000C00000000C",
INIT_02 => X"110400121014A411074204280042010000801104540220240024000080010042",
INIT_03 => X"40000888000041002040009302000181042000000000000A8080000000100000",
INIT_04 => X"0355134A4410692C60861400000010000008000080000B0100800582072A2001",
INIT_05 => X"0000400020000000320064000000000008000000000000022000000000000000",
INIT_06 => X"802050500000000100000400420000000029400000010200802D8000000400AC",
INIT_07 => X"8C0518832A800212449004200C200A20CA81008000000000010000000004AA00",
INIT_08 => X"0004050000000000040008080800801400000012002000000000000085030080",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE7394D4E04C1148010440605A158D94040",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C88A1F83F000020022002200020000000040004000000480012A000000000002",
INIT_01 => X"081025A00054C8C6940202C06F000801A50080B037810465AA0C60C00000008C",
INIT_02 => X"110400125014A4110746042880428100008411010603302100248000C0030106",
INIT_03 => X"4000018800010400044000DB822095C1142000002000102B8080000000100000",
INIT_04 => X"0F9B1B4E8208012E62940800020010000008808100000A4120000502072F8000",
INIT_05 => X"0040400260000001BA0374000000000808000000002100024000000000000000",
INIT_06 => X"81A078504000000180002502604008800029E01000000210802D8000000400EF",
INIT_07 => X"000400832F6000410692403298002000CBD90000000000A0012200000004AF80",
INIT_08 => X"0004070000001180040001000000000000000002400000000000000001806000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE701B2B18095005C029A93123518991024",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C6CC00100206811133331111580000000000010084084480A320000000100002",
INIT_01 => X"083425A020C40812840552811060DB28A10144A08801F060003809C014000C2C",
INIT_02 => X"114400321014A4110742042803520800408011054102201449240000D4210342",
INIT_03 => X"4800000800016D300048A0880020041014200001832C10A85080020000104400",
INIT_04 => X"ACE2ED56765C846DC75B56AAAA00109204480849C007540130A62A020480A800",
INIT_05 => X"410A401226C400218203048800321448480029091490400A60042D9091BE225A",
INIT_06 => X"7599005002184000A1002402434028800004001004000208800D8032810400E0",
INIT_07 => X"A515688080020959648240201830A2E02001820C20C4104A01030C2424820080",
INIT_08 => X"0004270091B0008034044140101044020004801A0052341A8D194C821101530A",
INIT_09 => X"0000000000000000005FFFFFFFFFFFF83800001EF9FE0F76FC3ED7DDE4E5F8C0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C088000001600222000000005A0000000040014000000480012A000000000002",
INIT_01 => X"08002500004408028400828000600000A10020A00000A060000000C00000000C",
INIT_02 => X"1084000000002411040204000042000000801100000220000028000081010002",
INIT_03 => X"4000000800000000004000800000000004200000000000000080000000108000",
INIT_04 => X"000D873106394000021014000200100000080000000000010000000204000000",
INIT_05 => X"0000400020000000000000000000000000000000000000020000000000000000",
INIT_06 => X"0000001000000000000004008000000000000000000002008008800000040000",
INIT_07 => X"0000008000000000048000200600000000010000000000000100000000000000",
INIT_08 => X"0000440000000000040000000000000000000002000000000000000001000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE07BF7F78E54CEFD36FAFD17FCFC7CF320",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08800000060022222222222000000000040000000000400010A000000000002",
INIT_01 => X"08002500004408028400028000000000A10000A000000060000800C00000000C",
INIT_02 => X"1004000000002411040204000042000000A01102160220000020000080010002",
INIT_03 => X"4000298800000000244008800000000004200000000000000080000000100000",
INIT_04 => X"0000008000042B24218800000200100000080000000001450000008A04000011",
INIT_05 => X"0000400020000000000000000000000000000000001000020000000000000000",
INIT_06 => X"0000001000000200002004000000000000000400000102008008800000040000",
INIT_07 => X"0000008000800000048000200000080000210000000000020100000000000000",
INIT_08 => X"0000040000001000040000000000000000000002000000000000000001000000",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"05104816EA00C199999999998B82D55555055577C0000675C3816AAAAAB80003",
INIT_01 => X"8014102000081213688B1862C400120ADA22C61962221218A90010E0957F0E0E",
INIT_02 => X"C200BAC50001061C8901300A2C0980A50085C801003641100400A00980206443",
INIT_03 => X"E2D5423CB284889002E20281C02900E8CC00000340A9401040162E6680824001",
INIT_04 => X"DAC651494D654F010FCA0208282AB2000D98181C14FDFC29876BFE33310017A2",
INIT_05 => X"0162E5846A0444221C5838881100401021048000000145D30AA9290000198B2F",
INIT_06 => X"84140A00A840000022800281241080040000104000002F219092A594094A9406",
INIT_07 => X"00000001010104011A42801D0244100440014000800490D0B58C444000A08004",
INIT_08 => X"612A8AB000AC00B4C66130400020000011002743150000000000100000548522",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE0334A4A0C60F6FB363875D4C538399B91",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4F74BF57E6E587FFFFFFFFFF92D71999998E665DC000E1D9E8758CCCCCF80000",
INIT_01 => X"2ADE30F033C915094A13393EDEF4B2265284CE4B6F40B85001AE0AB1FA003513",
INIT_02 => X"664123B786736A3991E3A47C1D59727F83855D59A1AC21CA6C30AAA2F8F149E3",
INIT_03 => X"01EF407061DE98DF4182021FC45117E22A0888D2C6F8E0FE6823B275CDE77725",
INIT_04 => X"D90A855E9396159B5AEBFD777C19EBC03DF139380EEDFC180363FE101FCE17A2",
INIT_05 => X"078D83F7F3CEFAFFFC5FFB96EBC021EE7D7ED00008BD6BB0067A7300009CCDED",
INIT_06 => X"5FEBF17BF430142FF1415AD12C11700001FFC007E7FAE8210DCA47FF1E58E6B8",
INIT_07 => X"105801B3FEE93C0112E1DACF82C6D945FFBB0E504085A1D076041DC000A6CE27",
INIT_08 => X"E66D1FC40024DFE9C023F3F007600088771815600D0020100800010630ECAF77",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE00C363180DDE2F82193AAC100343592A0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"80900040060040000000000040039E1E1E0F80060E1C067E2F81CF0F0F000003",
INIT_01 => X"82500F0000100211A6110064200002886984501A10005048A99041D0557F0A28",
INIT_02 => X"C0404B0000108804C04211220424A28000C0804940226454001080009001A502",
INIT_03 => X"6078001C3080000000EB02801129001CDC40000100810011D008380302004002",
INIT_04 => X"A662F955E7094500A5D54008A007F014021880C4040200098204001310000002",
INIT_05 => X"5062E0880ED505001C0038001036D20000002A1A1500108301F98CA1A12F1240",
INIT_06 => X"A4150A040AC0C8020A920A081014C00C2080386000000B2A5882A400218B3806",
INIT_07 => X"00500000008200051B06814AC10000000020810D82484020198561286D113146",
INIT_08 => X"266BAC10A190201046240000001405208005018303969048A41A4C084AD08000",
INIT_09 => X"0000000000000000005FFFFFFFFFFFE00917109AA06CA940889D014484C5D990",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"00014020080007FFFFFFFFFF82D7E01FE008005FC000E7E1C1F5F00FF0380003",
INIT_01 => X"0000000000000004108800000000000104220004006A80000000000000000000",
INIT_02 => X"00009440000005400C0000020400000000000000002200000020000940000000",
INIT_03 => X"6040001C3080000000E20280000900000C000000000000000014440010000010",
INIT_04 => X"018F03201F7C056400DE0C82A800700000180004040000098200001310000002",
INIT_05 => X"0000E08000000000000000000000000000000000000000830018000000302240",
INIT_06 => X"000000000000000000000100000000000000000000000B20831BA40000240100",
INIT_07 => X"0000000000000000000000100000000000000000000000001184000000000000",
INIT_08 => X"2110402000000000462000000000000000000103010000000000000000000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE02EDADE84C87AAA0501480081CC8CB890",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"00000000000007FFFFFFFFFF82D7FFE0000FF85FC000E7E1C1F5FFF000380003",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000027C00000180004400007E00000000000000000000",
INIT_03 => X"E7C6867DF780000093E60380000900000C000000000000000000000000000000",
INIT_04 => X"A01182938901EA66400042A800BFF000001800043F10023B8E18013770310046",
INIT_05 => X"0000EF8000000000000000090000043020040000000007CF1FF800000401401A",
INIT_06 => X"000000000000000000000000000000000000000000001F200002A40000000000",
INIT_07 => X"00000004012900000000000000001004004B400000101001F99C000000000000",
INIT_08 => X"E0040100040C4805EEE00000000000000000230F3F0000000000112000000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE0402621121D803000120200200848E033",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4410801502168D555555555520D7FFFFFF90001F8000057F8D55FFFFFFF00002",
INIT_01 => X"8880BE000439376128C090A2E09240284A30242970600098540084F0017FA04B",
INIT_02 => X"0511481A600817F8800B64437D11428202208800047EF900C80488000085480F",
INIT_03 => X"E7D80EFFF7CC20E513E60BF2044D11000C800040108C0022022B789ECAA60068",
INIT_04 => X"A339708A60102128A000100000BFF000281B33343C01007B8E02003FFA280436",
INIT_05 => X"0400FF909010C50924424A0A4E0001004202001000202BC71FF8010000B8224A",
INIT_06 => X"803440026C000403008142D00504C00C20E91842A2A29FA1D882B4013A0BC088",
INIT_07 => X"21004806380200410AC4DA18814000418A00800040002047F9DC000040152848",
INIT_08 => X"F7F9E20001A3C285CFE02200024000A2D500B307BF0020100800000000F05610",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE038888C1EF9FE0FF6FC3CD7FDFCFD78DB",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"6CD0E84501520D555555555524FFFFFFFF90009F8001C17F8055FFFFFFF00000",
INIT_01 => X"0A94BEAFE77D3C314A43D337A45241685290F4CFD22090F85C488C03D57FAC62",
INIT_02 => X"F6157F9A78589FFDD14B756901537001E028C4415900AB14E83DA22A50A5694B",
INIT_03 => X"0827A802001090086000807A1124150890A222023DA002AA52AE78DFEAF6314B",
INIT_04 => X"AFBB390A30488569A60142AAAA0003022943B3B043B10100111A80008AA81AC0",
INIT_05 => X"052A101242D56D8BA4574A886E20405943422101103308000007AC10111C264A",
INIT_06 => X"95B9400000680303A0700FD92A012001036D0602A2A68081D98111502ADFFEA8",
INIT_07 => X"84170066A882B0892642407D02A2B185AA202C00A20445CC006054040096280A",
INIT_08 => X"17FD23001023D3900105A3409342604044500400800084422111088C6164DF12",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE07B77739EF5EEFB76BAFF15E4BCFDF3A8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"8A99D0720284A800000000006A000000005FFF400C1804002D00000000000002",
INIT_01 => X"A00080000420E3E7BC8241B640909201EF20906F206006E5F4E2B4F0200040CD",
INIT_02 => X"A39050087D451C8190084003FC04B16802C11910167EDC8180382AA20006800C",
INIT_03 => X"E7C02FFFF780000017EE0BA0044D00122CC888D0700CC010020D0094F2A38B73",
INIT_04 => X"0CCAAD86201C00280300100000BFF010001A02043C0C517F8E6028BFF0000017",
INIT_05 => X"4000FFC89801B282044400068092100014108808048043C71FFF818080920000",
INIT_06 => X"41040000420040000B034B10850100000010002000013FA88082B4013ADFFF40",
INIT_07 => X"000000000008000109A00A58044208000002004400420003FDFD002024201006",
INIT_08 => X"E000800080100005CFE00000001004A091043B97FF1200000008000002F83400",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE00000000000000000000000000000001B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010800820001080000840037C00000000000000007E88008380000000040008",
INIT_03 => X"E7C0067FF780000013E603A0000D00000C800000100000000210008001000040",
INIT_04 => X"0065E581003800000200100000BFF000001A02043C00003B8E000037F0000006",
INIT_05 => X"0000FF8000000000000000000000000000000000000003C71FFF800000300000",
INIT_06 => X"000000000000000000000000000000000000000000001FA00262B40281000000",
INIT_07 => X"000000000000000000000002400000000000000000000001F9DC000000000000",
INIT_08 => X"E000400000000005CFE000000000002091002307BF0000000000000000000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE01D1A18B4B598CC60523ACB39BEBD603B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010000820001080000840037C00028600040000007E88008000000000040008",
INIT_03 => X"E7D8067FF7DC38FD53E623A0000D00000C800000100000000200008000000040",
INIT_04 => X"0000600C600421202100000000BFF000001A02043C00203B8E001037F0100426",
INIT_05 => X"0000FF8000000000000000191120214040200010000027D71FFF890105B40080",
INIT_06 => X"0000032FBC009428008000005014C00C2080184000001FA00002B40000000000",
INIT_07 => X"A5414910100200586004900081100AE00400800840802001F9DC000040010060",
INIT_08 => X"E002201C05A0000DCFE00000002000229108A327BF0230180C100C0000002200",
INIT_09 => X"0000000000000000003FFFFFFFFFFFE020272920E9ED0B200C52CF20B83A81DB",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"85F820440E61E5DDDDDDDDDD81D7FFFFFF8FFE3FDEBCEF7FDFD5FFFFFFF80007",
INIT_01 => X"AA5E3FF033CC1A1BA4993AAC8064328EE9265EAA400ABA7000401AC1DE00573E",
INIT_02 => X"F645FFF78F73EF7DDDE3B57E7C6F72BF89C15D49E0FE675E24302AA9F8D1E5E3",
INIT_03 => X"E7FFD67DF7DE1ADFDBEF578C5479263E7E600053CEFDE25C78BFFE7FDFF77F3F",
INIT_04 => X"F000600019C294D19C21E3FFFDFFFBDD7FF9393C3FF980BB8F5BC0777CC057EE",
INIT_05 => X"76AFEFFFBFDFFFFEC44D899FFFFFFFFE7D7EFEBEBFDE7FFF1FFBFFEBEFFFFFFF",
INIT_06 => X"1ECB83FFBFF5FD6EFED75ED91C9CF11D68861AE7475A7F2FDFDBE7EFBFFFFF30",
INIT_07 => X"525A85B4C00BBCA59DE7DBED41CEC5553003EF7FD6FFF159FF9DFDFAFFB34067",
INIT_08 => X"FFFFFFFDEFFFFFFFEEEFF3F2377C0F29F31F676F3F9DBA9D6EAEBF7E7B7C8F77",
INIT_09 => X"0000000000000000003FFFFFFFFFFFE0034B422CD53444E373420BBD2C2CFAB3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"11200008002844CCCCCCCCCC80D7FFFFFF8FFE1F5AB4AB7F5ED5FFFFFFEA8015",
INIT_01 => X"080A0E5012800008002029000029049200080A4000142822000002090A800110",
INIT_02 => X"4441D8370DC3416110A004547C8854AB88011100A0FC000A040022202A1000A0",
INIT_03 => X"97EF9671EFDC1ADDDB97570404512A062A000057CA7F0844783D024B19456E38",
INIT_04 => X"F000600019C294D19C21E3FFFDFFEEED6471292A3FB880BA4F598074784056EE",
INIT_05 => X"B08F8FF597FFB2B2410480BECEADCE767554B6B6BBCC7BEC9FFBBF6B6BFDFF7F",
INIT_06 => X"0E4383AFBDD5BD7A76D7C05C1CACF55C688218EC0C023C267842452AEBF3DE10",
INIT_07 => X"5A189424400B2A2290A9DE0561CCC5511002CAEB96BD5119FE1CEE9ADBF94076",
INIT_08 => X"FFFF31FD6BEFE677E8EF78FA3E4C8B1D1113474C3F2DAA956AA6BB7AD42E0FD3",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE03F1110E441278421012A097022228883",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4128400000606088888888888000000000000000420526004380000000080003",
INIT_01 => X"220A20501184080808802A90006000C202200AA40000A820004A02822A004110",
INIT_02 => X"B24427A5000A440440A21114001A00002288C440A980220A0CA1088828B120A2",
INIT_03 => X"0000000000008000800100041110020C8222220186D182D428827A14E2B25403",
INIT_04 => X"50000000098210901820A155540009C40D2018180000A0000001100000500000",
INIT_05 => X"15A5002D0D0A4D38405082013104A72722261202091E1438000012202401D9B5",
INIT_06 => X"0A46800000B00800500004000001100103520206A6A480028100406810240010",
INIT_07 => X"104A014050019880140100200006500414006601401B30140200388809005000",
INIT_08 => X"0000D0E0240C34682002D2B0852621C8444918E8000400400012112631000041",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE02064636888C821822C1405C480005B40",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A5F0A0540E75C5DDDDDDDDDD81000000000FFE20C60C677EC3D5FFFFFFD80003",
INIT_01 => X"805E1FFFF1C81619E659392E8076B2AE79965E4B402AB858000A0A71FF7FBF3B",
INIT_02 => X"E240FFF78F72EB588DE1A03E016D627D81408809E0FE455E66100001F850C5E1",
INIT_03 => X"E037C67C104E00C793E9038C403806345E4000438F5D604C281FFE7FDFA35F3F",
INIT_04 => X"F0000000098210901820A15554BFFBD43EB9191C03F1A03B811BD0370CD013C6",
INIT_05 => X"5285E07FAFDEDDF4C409891B75D6B6EE3D3C5A0A0D9C1FFF0003F2A0A4BFFBFF",
INIT_06 => X"1ACE817992B0592EDA015AC90010100001160005455A5F0B5E9BE3FFAE2BE130",
INIT_07 => X"100800B0D0011C0519C74BCC4004400034014755405DB059FF813DE82D92502F",
INIT_08 => X"17FFDFE8A4BFFFEDEE03D1B0173405A8A20D37EF00941008040A15263A748175",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE0F480845EF1DE1EFDF8B9DEFDFCFDF890",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000222222222225A00000000000140000000800020000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE03B7F7BFCFDFCEFE37F7E0FFDBCBDF3E0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"60008010001404444444444400D7FFFFFF8FFE1F0810817F0C55FFFFFFE00000",
INIT_01 => X"08800E0FC20105004A40000200128020129000010020000800000030017FA801",
INIT_02 => X"4401D8120D410161100004407D1050EB80011110017C00804A00222200200800",
INIT_03 => X"87EF8671E7DC18DD5386030004410002280888D2492C0080503D004B19452A38",
INIT_04 => X"A000600010408441840142AAA8BFE200205121203FB8003A0F588034780016E6",
INIT_05 => X"010A8FD092D5B2820004009ECEA040505450A01010806BC41FFBAD0101BC264A",
INIT_06 => X"0401032FBC40952822D340581C04E00C20C0186000003C2058420512ABD3DE00",
INIT_07 => X"00100004000A200000A0DA0541C081410002884882844109F81C440040B1006C",
INIT_08 => X"F7FF211C01A3C215C8E5204012400000111007043F00A05028100808402C0F12",
INIT_09 => X"0000000000000000001FFFFFFFFFFFE000000000000000000000000000000003",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


end;