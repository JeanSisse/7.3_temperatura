library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_master is
	port(clk             : in  std_logic;
        address_a       : in  std_logic_vector(31 downto 2);
        enable_a        : in  std_logic;
        wbe_a           : in  std_logic_vector(3 downto 0);
        data_write_a    : in  std_logic_vector(31 downto 0);
        data_read_a     : out std_logic_vector(31 downto 0);

        address_b       : in  std_logic_vector(31 downto 2);
        enable_b        : in  std_logic;
        wbe_b           : in  std_logic_vector(3 downto 0);
        data_write_b    : in  std_logic_vector(31 downto 0);
        data_read_b     : out std_logic_vector(31 downto 0));
end; --entity ram     

architecture ram_master of ram_master is
signal enable_a_lo       : std_logic;
signal wbe_a_lo          : std_logic_vector(3 downto 0);
signal data_write_a_lo   : std_logic_vector(31 downto 0);
signal data_read_a_lo    : std_logic_vector(31 downto 0);
signal enable_b_lo       : std_logic;
signal wbe_b_lo          : std_logic_vector(3 downto 0);
signal data_read_b_lo    : std_logic_vector(31 downto 0);
signal enable_a_hi       : std_logic;
signal wbe_a_hi          : std_logic_vector(3 downto 0);
signal data_read_a_hi   : std_logic_vector(31 downto 0);
signal enable_b_hi       : std_logic;
signal wbe_b_hi          : std_logic_vector(3 downto 0);
signal data_read_b_hi    : std_logic_vector(31 downto 0);
signal address_a_reg     : std_logic_vector(31 downto 2);
signal address_b_reg     : std_logic_vector(31 downto 2);
signal enable_a_lo_256       : std_logic;
signal wbe_a_lo_256          : std_logic_vector(3 downto 0);
signal data_write_a_lo_256   : std_logic_vector(31 downto 0);
signal data_read_a_lo_256    : std_logic_vector(31 downto 0);
signal enable_b_lo_256       : std_logic;
signal wbe_b_lo_256          : std_logic_vector(3 downto 0);
signal data_read_b_lo_256    : std_logic_vector(31 downto 0);
signal enable_a_hi_256       : std_logic;
signal wbe_a_hi_256          : std_logic_vector(3 downto 0);
signal data_read_a_hi_256   : std_logic_vector(31 downto 0);
signal enable_b_hi_256       : std_logic;
signal wbe_b_hi_256          : std_logic_vector(3 downto 0);
signal data_read_b_hi_256    : std_logic_vector(31 downto 0);
begin
process(clk)
begin
if rising_edge(clk) then
	address_a_reg <= address_a;
	address_b_reg <= address_b;
	end if;
end process;
data_read_a <= data_read_a_lo when (address_a_reg < x"0001000"&"00") else
data_read_a_hi when ((address_a_reg >= x"0001000"&"00") and (address_a_reg < x"0002000"&"00")) else 
data_read_a_lo_256 when ((address_a_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_a_hi_256 when ((address_a_reg >= x"0003000"&"00") and (address_a_reg < x"0004000"&"00"));
data_read_b <= data_read_b_lo when (address_b_reg < x"0001000"&"00") else
data_read_b_hi when ((address_b_reg >= x"0001000"&"00") and (address_b_reg < x"0002000"&"00")) else
data_read_b_lo_256 when ((address_b_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_b_hi_256 when ((address_b_reg >= x"0003000"&"00") and (address_b_reg< x"0004000"&"00"));
enable_a_lo <= enable_a when (address_a < x"0001000"&"00") else '0';
enable_b_lo <= enable_b when (address_b < x"0001000"&"00") else '0';
enable_a_hi <= enable_a when ((address_a >= x"0001000"&"00") and (address_a < x"0002000"&"00")) else '0';
enable_b_hi <= enable_b when ((address_b >= x"0001000"&"00") and (address_b < x"0002000"&"00")) else '0';
enable_a_lo_256 <= enable_a when ((address_a >= x"0002000"&"00") and (address_a < x"0003000"&"00")) else '0';
enable_b_lo_256 <= enable_b when ((address_b >= x"0002000"&"00") and (address_b < x"0003000"&"00")) else '0';
enable_a_hi_256 <= enable_a when ((address_a >= x"0003000"&"00") and (address_a < x"0004000"&"00")) else '0';
enable_b_hi_256 <= enable_b when ((address_b >= x"0003000"&"00") and (address_b < x"0004000"&"00")) else '0';
wbe_a_lo <= wbe_a when  enable_a_lo='1' else x"0";
wbe_a_hi <= wbe_a when  enable_a_hi='1' else x"0";
wbe_b_lo <= wbe_b when  enable_b_lo='1' else x"0";
wbe_b_hi <= wbe_b when  enable_b_hi='1' else x"0";
wbe_a_lo_256 <= wbe_a when  enable_a_lo_256='1' else x"0";
wbe_a_hi_256 <= wbe_a when  enable_a_hi_256='1' else x"0";
wbe_b_lo_256 <= wbe_b when  enable_b_lo_256='1' else x"0";
wbe_b_hi_256 <= wbe_b when  enable_b_hi_256='1' else x"0";



ram_bit_0_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"88280C4C7B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"00160090920C04800904848262220277E05152B280780D407428E723C01E1400",
INIT_05 => X"0006D46207801E400183C0707800E6000E008057641E00473C40680D32330C00",
INIT_06 => X"203F70C165000225E2C11E2C12A0D0144AC27206582C166504800000B0FC21D5",
INIT_07 => X"920CFC5E6D233B964E7CD99DFB870E1DDDD889C5FBDC440129A0604442180238",
INIT_08 => X"80B036AD23C17544C581000657A0E8E83D86F0E4A7B2D88AAAFD7FE0E1833AC5",
INIT_09 => X"C800016D82082E2081B6C0027ADA398000008A504318404005B70663212C04A0",
INIT_0A => X"4AF4AA414568729139FAD610C00001A2502440888420247041E87681008CE9AF",
INIT_0B => X"00890022B826E250B12346F1244812240912048941621804A150CA1CA45C254D",
INIT_0C => X"B2E0F1F80FA97FE0F0009E0FC40FA97FE0F0009E0FC048211E9C11C31F82E4A0",
INIT_0D => X"C3CB5F040FAB3FE0F0009E0FC40FAB3FE0F0009E0FCC42EFDFBF0AE03080E2AE",
INIT_0E => X"187806013879BA878FE807F65FBF12E0380231F0BD9E3FC08FEBD6F661C0E008",
INIT_0F => X"C83136B248831ACBFC8BBDCAB779BC699F20180309A0F83BE2B87C7C42EFDFBF",
INIT_10 => X"9947184131B59003FFEC07F00003F01FB90BE9F01FC8B38C2098DAE007F323A0",
INIT_11 => X"D065703080E29F1B2BE9F8A27E6E915C0E004C72BEC800FE7464290626D7003F",
INIT_12 => X"6F846DFC0C2352A0024B83F07F198BE9F8A0FFDA2A3C0202B8776A2FA7F023F7",
INIT_13 => X"11800014481A6105810941C5C068000CD4004C0905E52630BB1AE49C2BA7F98D",
INIT_14 => X"7E96656074EA560F0416A24844B01302A26100C4801844069B0C88881A28C141",
INIT_15 => X"E2781EA781E2781EA781E2781C33C0613C0E21020800239450116ED443C041B4",
INIT_16 => X"8112C1241140A056954AB0C280D0002020187007122C3E04E03383E2781EA781",
INIT_17 => X"1204812048120481204812048120481204812048120481204812048120481205",
INIT_18 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_19 => X"4000000000000000001204812048120481204812048120481204812048120481",
INIT_1A => X"10410411062084E57CE2641DC71C71574E09B56C74DAB16782171CF13043A85D",
INIT_1B => X"F87C3E1F0F87C3E1F04104104104104104104104104104104104104104104104",
INIT_1C => X"0007C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0",
INIT_1D => X"0000000000000000000000000187C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE500",
INIT_1E => X"BD54BAF7FFD55EF007FD75EFFFAE97555557BD75EF5D00000000000000000000",
INIT_1F => X"FFC0000AA843FE00AAFBE8B45AA803DFEFA28428B455D0017410A28428AAAA2F",
INIT_20 => X"57FFFEBAA2D5401450051401555D7FC0145F7AEBFFFF08002AA10A2AABFEAAA2",
INIT_21 => X"5D7BD755555517FFEFA280021FF082E974AA5D7BFFE000804000BAAAAAAAB455",
INIT_22 => X"A5D2EA8B45005168A10AA8028A10087FD7410557FC21555D51574AAA2FFE8B45",
INIT_23 => X"FFFFAE95410AA80000005D003FEAAFFAEBFE00A2803FEBA002A820AA0800174B",
INIT_24 => X"5EFA2AEA8A10000417410A2FFE8BEFF7FFE8B45FFFBC00005D003FF45557FC01",
INIT_25 => X"000000000000000000000000000000000000000000557DF5500003DFEFFF8417",
INIT_26 => X"12555F524AFE38B780154BAFFF1D54AF0075D75EFEBAE9554540754717F1F800",
INIT_27 => X"B6AB50B6AABDE12BEA0AF010B7D1F8F47E00A2DB45AA8A3AFD7B68E2AB78550E",
INIT_28 => X"A43FE9257F1E816D557095EAAA2D1401D500002A150038038E285D7F78FD7000",
INIT_29 => X"57545A87AAD178A8002D1D21C5E8257D5C7AA854008700249243A412EBFF5542",
INIT_2A => X"02D152A82000E3A5D2150AB8F401471EDBC0B680900AAF52B474385D75C502D1",
INIT_2B => X"D417FD7E9541242FE920AD082E10A28F6A150012A2F02AFFDF40E85F475451D5",
INIT_2C => X"55080550E87B7A405B52AAD152BD00151EAFEDB52E3F1EFFFF485A2DA3D5D24B",
INIT_2D => X"445057F40545850000000000000000000000000000000000000000000005AAF5",
INIT_2E => X"AB55F7AEAABFF5D2A81151FB8635A02FA69574BAF7D5555AF0D79D55FFA2AC97",
INIT_2F => X"34A08D46F6ABE7082AAAAF2FAC77FE00FF16565B2FA9075F4F7B3EBDF50FEAEA",
INIT_30 => X"C95256803CE3AEB038662E5D81406014D5D51F5E08A394003A908B8410E707EF",
INIT_31 => X"C0954AF0151555AF58794040077D774FAE8C798A11A0EAEF75F7AA84001A7052",
INIT_32 => X"245B4E1870108B11020AD4AA05542A0A05051023F9A9D57B63BFBF906CB45FAB",
INIT_33 => X"ABD5F5F0DA6BC9525688C1A2A0C06E9FEE5555BE48AB2A2AE0A0F20C43EAC562",
INIT_34 => X"0FF8000000FF80F55E25C00A0BA7FBED407A97F6F35F498B96BEB12DAAB77558",
INIT_35 => X"00FF8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF800000",
INIT_36 => X"000000000000000000000000000000FF8000000FF8000000FF8000000FF80000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000800000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"CA1800080848B0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000010822C00803804000001999EF9C00040B0002000001000640200001018",
INIT_05 => X"0000400244000000014200004000000004000000001000032000200002100800",
INIT_06 => X"202800208500000080412804100CB08000302220080408010000000404100844",
INIT_07 => X"25FC4C5AF6FEF002230018010860C1833C460044204C000008A0041000080008",
INIT_08 => X"0010008D22C0F55000010000524481890BC000263000188AAAA10F8C1830562B",
INIT_09 => X"041001B102002E20013600022D8819000000A000110A4000002C204000240420",
INIT_0A => X"0BE0B002605C1C1108484400C000002040040820000020104100028800002801",
INIT_0B => X"000000081001004010810510040802040102008100200800A1100707040101E2",
INIT_0C => X"10F18058000003C0F000A000C4000003C0F000A000C0000012187087010AE4B0",
INIT_0D => X"00012704000003C0F000A000C4000003C0F000A000CC4200002F08E030800000",
INIT_0E => X"1878060000000AAC00680000001F10E038000000078808C00000023461C0E000",
INIT_0F => X"4800025200040A00D000000202090C281F201803000000240218C0044200001E",
INIT_10 => X"904618400012900001EC03F000000000392100B00048230C200009A000130320",
INIT_11 => X"806070308000000961002880204A901C0E00000002C9000260640900004D0000",
INIT_12 => X"0904285C0C0312A002000000083881002880025A0A3C020000002A8400B00007",
INIT_13 => X"08400004080030008010468220A00008D0000801046004308A18500002012800",
INIT_14 => X"2200000840280206089000004090110200000000001454000200828008081110",
INIT_15 => X"A4191A4191AC191AC191A4191A00C8560C8D2910000060901010401E13405111",
INIT_16 => X"8000410410028000100800140000002004103224002006406401918C191AC191",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"0000000000000000000200802008020080200802008020080200802008020080",
INIT_1A => X"1451455901218D2C4CA2900C9249258306BABEFC54A081701C397452B4008A04",
INIT_1B => X"BADD6EB75BADD6EB755555555555555555555555555555555555555545145145",
INIT_1C => X"0005D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2EB75",
INIT_1D => X"0000000000000000000000000607FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF600",
INIT_1E => X"E80010AAAABFFFFFF803FE10F7D17FEBA55556AAAAAA80000000000000000000",
INIT_1F => X"2EBFEBAFFD555400557BD54BA5D7FFDF45A2FBD75EFA2AE97555F7FBFFF45FFA",
INIT_20 => X"A802ABEFA2D568A005D5157400AA8028AAAF7FBD54AA002A955555D7FE8ABA08",
INIT_21 => X"FFFFFDF55AAFBC0010555540010550417555AA8028BEFAAAE97555082A80000A",
INIT_22 => X"A557BD7410550428ABA5D5168ABA552EBDFEF5D7FEAA00AAAABFEAA007BC0145",
INIT_23 => X"FFFFFFEAB55557FFFEBAAAD568B45A2D5575555D7FC2155F7AEA8BEFAAAA954B",
INIT_24 => X"4AA5D7BD74000804154BA082ABFF55FFD57DF45F7D568ABAF7AABFFFF082ABFF",
INIT_25 => X"0000000000000000000000000000000000000000002EBFFEFA280021FF082E97",
INIT_26 => X"95545E175EFF57BF8FC2000BEA4BAE97F78A3FE28E3D17DEAA485FE8E02B5000",
INIT_27 => X"FD55455571E8A2A087BF8EAAEB8E0016D5D75D54BA5D7BFFF7DA2FFD55EFAAA4",
INIT_28 => X"AA07157428145A00AA8A2FBD7B6DF6AA28550E10405F7A4AFE38EAA0924921C2",
INIT_29 => X"6AAB8E971471C7010B7D168F47400A07A28415A001684104155C5B6DF6DBEFBF",
INIT_2A => X"5FD4BFBD7B6A0BF492415FC20105D24AAABF1FFBC7010FF8A38FEF557FEAB78B",
INIT_2B => X"FE38017EBA4A8EB8F6FFD5FE8B7D557495EAAA2D16D1FDBED56A55557A43DE38",
INIT_2C => X"C7AA854008700249243A417FFF41542F5D717FE2AAAA56DEBD17FE3DF7FB7FEB",
INIT_2D => X"FBA007DFCA127B8000000000000000000000000000000000000000000002A3D5",
INIT_2E => X"FFEFAAFBD55FFAA8416545A6FB60F47AF2A00010F78028B15F7823FEAAA2D57D",
INIT_2F => X"21A022A38C20B2552E975F758516AAAA0869AAAB8A7C19C55550E8574BA557BF",
INIT_30 => X"895755FFEFBCEE5FBAACB10085EE5DE10A2AEBFF55F7BAAA8565DBAC1112FFAC",
INIT_31 => X"02EABEA097BEAAFAF2863FA00DD574201E7AD1FFF5575841DE08007FC2048002",
INIT_32 => X"AF9554FF57EFBFA18D4FBFFF40FF809D4000D7FC00FC5D062BBA05ED5034472A",
INIT_33 => X"FED17DFBFF6963FCAAA2283CF14050062B0A2F7AE8B5D5D51F5E18ABD5EAFFF2",
INIT_34 => X"0000000000002CB75F7AA84001A7052C95256807DC31AA8114DE55F5BED201FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000800000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2812",
INIT_01 => X"0005A18A0849204D1CA024A542500368404000720885800802000106E4D10204",
INIT_02 => X"5C010802020408040C600850AA055254090541A111240A104A0000000908B510",
INIT_03 => X"182202210800004401060A0010041028021560A0218808002440840008C80550",
INIT_04 => X"21030A008814500120A06B0870201010258261E141A2326511024182142494D2",
INIT_05 => X"48484098142953388552102442884882B58A09291290A1120A81A3C200418DCA",
INIT_06 => X"22208802800554529001C9003A2800203120000104810100002A614008102244",
INIT_07 => X"0008040000221040408100890C0000011804480420420154000088096A0EA8C0",
INIT_08 => X"B846C0081190C105424705510A08828A0B190C0428040080A0A10F8000009200",
INIT_09 => X"20B0573165541CD54822160A89E89020AA8A80CA9D39CE215264B15818004442",
INIT_0A => X"0402100C088104010AC80005C568147007031012D40D71824114081538000048",
INIT_0B => X"550055481205100C000134128304408020C11020040244D00001306100A24600",
INIT_0C => X"00500000B01480010000A00001501480010000A0000801487334E34C1A980001",
INIT_0D => X"00012001501480010000A00000B01480010000A0000138000040000800000000",
INIT_0E => X"02000000000000A00003600180400010000000000608000A5004090008000000",
INIT_0F => X"000002400008C4000220420040800280001000000000002400000001A1000040",
INIT_10 => X"2090000000120C94000200000000000001380001C01048000000090298040440",
INIT_11 => X"2018000000000001580002508010440000000000000953008088000000481380",
INIT_12 => X"10180000820080000000000008201800024C000100000000000002E000095000",
INIT_13 => X"09130A82000C90A0000081A004342AB001720040000000000001502050000422",
INIT_14 => X"094882958000934200904407600090822085E0100D52498002B1041092001514",
INIT_15 => X"3C1011C1013C1011C10134101140801A0808AD4451394CD0391A541593C04B59",
INIT_16 => X"022810800000A0289A6D084D4021208106142034406144004041011410114101",
INIT_17 => X"4010040104411044110441100401004010040104411044110441100401004010",
INIT_18 => X"0102401024010241106411064110640102401024010441104411044110040100",
INIT_19 => X"2F81F81F83F03F03F04110641106411064010240102401024110641106411064",
INIT_1A => X"0820823047486021658010816596597700138D70C030B542923650C7D0002281",
INIT_1B => X"944A25128944A251282082082082082082082082082082082082082082082082",
INIT_1C => X"F804A25128944A25128944A25128944A25128944A25128944A25128944A25128",
INIT_1D => X"0000000000000000000000000787C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF871",
INIT_1E => X"5420AAAA843DFFFAAD1554005D7FD74AA0004001550000000000000000000000",
INIT_1F => X"2EBFF45AAAAA8A10A2AE80010A2AA975FF5D003FE10F7D17FEBAF7D5420AA085",
INIT_20 => X"D7FFFF45A2AA975EFA2FFD7555FFFBFFF45AAFBC20AAF7D1575EF55517DF555D",
INIT_21 => X"AAAE95555552E974105D517DF55AAAAAABEFAAD1575EFAAAE974AA5D51554BA5",
INIT_22 => X"F552E82010F7AABFE10FFD542145FFD5554AA555555555557FE8ABA082EBFFFF",
INIT_23 => X"EFF7FBC0010AA802ABEFAAD540000FFD540000AA802AABAF7FFC2010AAAE821E",
INIT_24 => X"555AA8028BEFAAAE821550851420AA002E800AA08042AB45007FC00BAFFD168B",
INIT_25 => X"0000000000000000000000000000000000000000002E80010555540010550417",
INIT_26 => X"7DEAAE95F40002157F470AABE803AE97A2DF55400557FD54AA1D04001C515000",
INIT_27 => X"E105EF55517DFC5552ABDF45B6AEAFFD5F7A482000BEAE905C755003FE28E3D1",
INIT_28 => X"A4070BA5FD0154BA5D7BFAF7DA2AE955EFAAA495545E3F5EFF57F7FE80082FFD",
INIT_29 => X"571E8AAF082AB8EAAEB8E0016D5D2A924105D5B7FF7DB6AAAABC7BEDB505EFBE",
INIT_2A => X"E80495038AAAEAF1D7410E80000FF8438E00B6DF68FEF4871D24BA495B5556D5",
INIT_2B => X"80071ED1EFEAF1EFFFDEAD1C5010AA8E2FBD7B6DF47A00EBDB50000A380AAE28",
INIT_2C => X"28415A001684104155C5B68E2DBEFBFFBC703AE2DF42AAA002A851C214003FF6",
INIT_2D => X"4AA550002155510000000000000000000000000000000000000000000002087A",
INIT_2E => X"215555003FEAAAAD57DEBAA2FDDC01051FBD74BAF7802AB05AAFBD5400557BD5",
INIT_2F => X"60F47AF7FC20B2F7FBC015D58517FF555D2ABDF55F782BEB47AFAD00010F7AA8",
INIT_30 => X"22A955FFFFC20FFF3AE544108410174BA557BEABEFAAEBD55FFAA1456547A2D3",
INIT_31 => X"D4420BA547FD75FF58516AAAA0828AAAB4A78016545540400010557BFDFFFF78",
INIT_32 => X"FFBD550AAFACAAA122AA8954BAA2AE9D545002A800A8FF862BA00F2F9E8F0050",
INIT_33 => X"002E954505C417FFFF08555555BAAD335B57AB5155400A2AEBFF45FFFB404007",
INIT_34 => X"000000000000061DE08007FC2048002895755FFAEBCFE57BBA57002DF3C4AAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000001000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B815602110494074133520400E02B92206",
INIT_01 => X"014C9BC048800168240442C99E004B61404040028804A0080A000516A0990A08",
INIT_02 => X"4809A900031800444440589866E331352180D468B8000E600C0081110B802CD0",
INIT_03 => X"DA16C0200C0001423583480408D60520320066810A80881068A808029C856330",
INIT_04 => X"2088681DA82740EC92307364B37569100A84E1E11C251210990040420E005A48",
INIT_05 => X"2D284A102414411A314A0A02C18C01B9854368280A506902018C2442484038D1",
INIT_06 => X"23600016801CCCAA9061C9061C0D0080001005210C8761001166CCC40C110826",
INIT_07 => X"0178045800B6540063000889082040A13A0716042440833280038C89904E6400",
INIT_08 => X"D20A480810804451421D1CC8024481994B5500061000088000A10F840854973A",
INIT_09 => X"2079CCB035E03CCC5D2A35620988100A698761C0953B6E84C82C404018304D42",
INIT_0A => X"070070202A90340440C80004CCE4CC1042061913208CE8024380880820010040",
INIT_0B => X"3302CCC01300104018900402870C4287214210E114200410EC20242D01015E84",
INIT_0C => X"4801000180148000000800100040148000000800100401C33249049051218073",
INIT_0D => X"04008001001480000008001000E014800000080010001C000040000000000000",
INIT_0E => X"0000000000004408000068018040000000000001400800091004090000000000",
INIT_0F => X"00004100812644000004400140800280000000000002000008008000B0000040",
INIT_10 => X"20900000020800CC0002000000000020400800030010480000010400C8040440",
INIT_11 => X"2018000000000060080004418010440000000000410015008088000008200540",
INIT_12 => X"80188000820080000000000100400800041C0001000000000000902000014C00",
INIT_13 => X"284B264208448260E27285A23224E660084208410000004444000E0000000020",
INIT_14 => X"0840024D810283021280400720C0348002854C001CC3158026A2040028090441",
INIT_15 => X"80901A0901A09018090188901A248054480C0C0041116DD0115E011599641E59",
INIT_16 => X"C6C8408514028028D06C0C5D20030BA1010021B000020402400501A090180901",
INIT_17 => X"4290C4290843908439084390843908439084390C4290C4290C4290C4290C4690",
INIT_18 => X"290C4210E4290C4310A439084310A439084310A4390C4290C4290C4290C4290C",
INIT_19 => X"5D54AAB556AA9556AAC310A439084310A439084310A439084210E4290C4210E4",
INIT_1A => X"0820825103A1600054C0F4012492490300C78C706428A1411133586294020A90",
INIT_1B => X"D4EA753A9D4EA753A92492492492492492492492492492492492492482082082",
INIT_1C => X"8086A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A353A9",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE024",
INIT_1E => X"5421EFAAFFD54AAF7D168B45AAAABDF5500002AA100000000000000000000000",
INIT_1F => X"043DF45FFD168AAA0855420AAAA843DFFFAAD1554005D7FD74AAA28400155005",
INIT_20 => X"2AA955FF5D003FE10F7803FEBAFFD5420AA080400155AAD5554AAF7802AB4500",
INIT_21 => X"AA8028B45A2AE82155A2FBFFEBA0800021550855555FFAA84001FFAAAE80010A",
INIT_22 => X"0085168ABAFFFBD54BAAAAE97400A2FBC20AAA284175EF55517DF555D2EBFE00",
INIT_23 => X"55AAAA954AA5D7FFFF45AAAA975EF007BD7555FFFBFDF55AAFBD55EF5D2EBFE1",
INIT_24 => X"BEFAAD1575EFAAAE974AA5D00175555D0015410F7AAAAAAA55043DE00FFFFD55",
INIT_25 => X"00000000000000000000000000000000000000000004174105D517DF55AAAAAA",
INIT_26 => X"D54AABC04001C51551471D7AAF1D05D2EBD56DB7DBEAEBFF551C042AA101D000",
INIT_27 => X"B50492EB842FB5508043FF55EBD56ABD75D5B470AABE8A3AFD7A2DF55400557F",
INIT_28 => X"8E82557FD2082000BEAE905C755003FE28E3D17DEAAEBDF40002550F47155AAD",
INIT_29 => X"5517DF40552ABDF45B6AEAFFD5F7A48017DAAFFFAE821C0A0717D1C5B575FFB6",
INIT_2A => X"F7D5C55D7492E90E3808756DA92EBFFD74BAE3AE85480FFFFC00AABE8E105C75",
INIT_2B => X"241043AE10EAF5C5547FF80954AA5D7FFAF7DA2AE905EF0075D5545E3F5EFF57",
INIT_2C => X"105D5B7FF7DB6AAAABC7BEDB505EFBEF5C7092FF801756D490A10438EBA4B8E9",
INIT_2D => X"F555D0028A00510000000000000000000000000000000000000000000000E124",
INIT_2E => X"8B45AAFBD54005D7BD54AAF78002155515157555AAD142040A2D57FFFFFFAEBF",
INIT_2F => X"DC01051AE955F7AAFBC0000AF843FF5500003FF55AAFD6AB455157D74BAF7AAA",
INIT_30 => X"E955FF557BD74EFFBACD41577B8400010F7AA8215555003FEAAAAC53DEB8A2FD",
INIT_31 => X"FEC20BAF7AA8015558517FF555D2ABDF51F782BCB47ABAE801FFAAFBEAA105D2",
INIT_32 => X"8554214FA2D3EAF57AFFDD7555082AA0AAA00557FEA8A2FDD64BAAF8282012AF",
INIT_33 => X"082A820AAAB842AA00000028AB0AAFF48547AE04174BA557BEABEFA2AA951FF8",
INIT_34 => X"0000000000002A80010557BFDFFFF7822A955FFFFC21FFF3BE40412DE02955FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000800000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303000048B3532C82D04A16002",
INIT_01 => X"210399800808004C1C20650E1E104368403008418984014902030006A8910200",
INIT_02 => X"480108A200000000444148E41E80F00A4104311868200200080000000988A390",
INIT_03 => X"0CA08220080000D004260A0240109028270012603000000030808C4208C000F0",
INIT_04 => X"4403A609A055306BC2C0735810CEE5100A0A48E16B8370E3808241D03845D002",
INIT_05 => X"ECE8698800791403AD3038AE079059A790E245A19A41E4120BAB86C00001D312",
INIT_06 => X"23208806000C3D220023C0021A21008891048C00040341121661E3C10000A064",
INIT_07 => X"0008045000220440000000090800102118400204A04100F040018019004B8001",
INIT_08 => X"0E11400810906441123323C0424190880B0108002000000880810F9002041200",
INIT_09 => X"22003C2309671584786E0F5A88889031EF9F05D884794FA03A24781810106D02",
INIT_0A => X"0409400E4282A00142400004DC3C82400702003200872003FB14080828400010",
INIT_0B => X"F050C3C00095000C008135040002010100800040001400C00401208800F01A14",
INIT_0C => X"08000002E0100000000800000220100000000800000001C87261C51C42390240",
INIT_0D => X"0400000280100000000800000360100000000800000035100040000000000000",
INIT_0E => X"00000000000004000000D8008000000000000001000000155000080000000000",
INIT_0F => X"000040000120EC00004002214000008000000000000200000000000094100040",
INIT_10 => X"001000000200050C000200000000000040080005800008000001000168000040",
INIT_11 => X"000800000000004008000448000040000000000001003C000008000008000D00",
INIT_12 => X"800800000000800000000001000008000017000100000000000010200002C800",
INIT_13 => X"150F5E0400101000227200800E271E00288400800208004C04C0080000000052",
INIT_14 => X"818082450000920280C544310041B408880EC51060461589225100063E9012D6",
INIT_15 => X"1410C3410C1410C1410C3410C100869A08618C00772201D899BA003591510A59",
INIT_16 => X"44E0110004480020986D4815044369A00006203041C3443043010C5410C3410C",
INIT_17 => X"0080001002008040100200800000060180000006008000100600804000020180",
INIT_18 => X"0000010060080201800000040100201802008040100201804000020180001006",
INIT_19 => X"64B261934D964C32698080401000000060080601800000040000201806008000",
INIT_1A => X"1451457A604C8D0C28A280CD145144C1863807E0500014385DAF345041488280",
INIT_1B => X"1A8D46A351A8D46A355555555555555555555555555555555555555545145145",
INIT_1C => X"1F60D068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D06A35",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE077",
INIT_1E => X"02ABFF087FFDF5508003FEBA087FD54BAAA84154005500000000000000000000",
INIT_1F => X"2EBFF5500003DF455555421EFAAFFD54AAF7D168B45AAAABDF55A2802AA10000",
INIT_20 => X"A843DFFFAAD1554005D7FD74AAAA840015500002AABA082E954005500021FF5D",
INIT_21 => X"FFD168BEF080028BFF0855555455500174BAA2AABDE0055517FF555555420AAA",
INIT_22 => X"0085168ABA0055574BA5555554BA5D0400155AAD1554AAF7802AB4500043DF45",
INIT_23 => X"AA5D0400010A2AA955FF55003FE10F7803FEBAFFD5420BA085168A00007BFDE1",
INIT_24 => X"1550855555FFAA84001FFAAFBEAB45002A97545F7D1555EF55043DF5555517DE",
INIT_25 => X"0000000000000000000000000000000000000000002A82155A2FBFFEBA080002",
INIT_26 => X"BFF55BC042AA101D0A28BC7007FFDF45080A3AEAA007BD2482BE84124285C000",
INIT_27 => X"4974004100021FF492AB8F7D1C0438E381451471D7AAFBD0492EBD56DB7DBEAE",
INIT_28 => X"557AFED1C5F470AABE8A3AFD7A2DF55400557FD54AABE84001C5550A28ABA142",
INIT_29 => X"B842FB5508043FF55EBD56ABD75D0428BEF005557545490012482B6A0BAE2849",
INIT_2A => X"557F6DA101475FDE10145F68A921C55504924955524AA140E0717DAADB50492E",
INIT_2B => X"F5D043AF6D405F78E3A1C2002000BEAA905C755003FE28E3803DEAAEBDF40002",
INIT_2C => X"7DAAFFFAE821C0A0717D1C5B575FFB6DF425575D7BEFB55002097555FFD5401E",
INIT_2D => X"010F784000AA5900000000000000000000000000000000000000000000020801",
INIT_2E => X"2000A2D57FFFFF7AEBFF55FF8028A00512EAAB45007FFFF55082EA8AAA087FC2",
INIT_2F => X"02155512AAAA085D04174100800021FF002EA8BEF5D0428ABA595557555AAFBC",
INIT_30 => X"402000FF802ABAA04552ABFF597FD74BAF7AAA8B45AAFBD54005D7BD54AAF780",
INIT_31 => X"2F955FFAAFBC0000AF843FF5500003FF55AAFD6AB4551002ABEF005555555000",
INIT_32 => X"A843DEB0A2FD5600051537DE005D557DE005D7BE8AA85555400100879560AA59",
INIT_33 => X"000417545FFD5421FF5D0428BEF0079FCABA598400010F7AA8215555003FEAAA",
INIT_34 => X"00000000000004001FFAAFBEAA105D2E955FF557BD75EFFBBCD415521FBFDF45",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000001000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB0A0791B1B41694368283C81F9996A091A32152007AB37B20E07C0C1E002",
INIT_01 => X"881FBC449030884C446A00000034824841280A00084000C8C212812EEA953231",
INIT_02 => X"C809AD5CB118E640A4F408FC011FF0002080000082CCC66609DB7DDDCB1F2036",
INIT_03 => X"4A100E4D3E4C90D290831C824A4204720B20048A88800000B8E0F91028C5500E",
INIT_04 => X"00144884922644001914830051110A71E03040F0105B001C662AE22DC08A3408",
INIT_05 => X"120340220B88820041CDC451B860A6506BEBD08265AE105714505F0152122449",
INIT_06 => X"207F7890752C037372A1D72A398CD084C890EA2950A37E270660182C0D2C8080",
INIT_07 => X"9378355E64B66F96231CC81D2DAB468D38C601C5FFF54FF1C9A46490261C4B39",
INIT_08 => X"7F105CAD1089654115814FC60284A1A93B46F4621030C800001D7FA56891162E",
INIT_09 => X"E00A003C832D25328526C082DF9AB88C104024C09639441807B78661090C24A1",
INIT_0A => X"4FD32A2E2A9992944AF2D611C3FC01B2152109204C28B67061EC928920C569E7",
INIT_0B => X"F0313FE92C22F21CA0B363C0A242502028901408154218144D712664A5F15AC1",
INIT_0C => X"B2F0F1E01BE53FE1F000BE0FC41BE53FE1F000BE0FC80020130841840308653F",
INIT_0D => X"C3CB7F041BE1BFE1F000BE0FC41BE1BFE1F000BE0FCD806FFFAF0AE83080E2AE",
INIT_0E => X"1A7806013879BAA78FC103FF5F1F12F0380231F0BF9E3F02A7FFD63669C0E008",
INIT_0F => X"483136F200A822CBACAB9DDEB7F9BC291F30180309A0F83FE2B87C7D006FFF9F",
INIT_10 => X"D1C6184131B7980DFFFC03F00003F01FB931E9C1DBF8A30C2098DBE2FF7F2320",
INIT_11 => X"F060703080E29F1B71E9F6427EFE901C0E004C72BEC95FEF64E4090626DF15B7",
INIT_12 => X"EFAC6DFC8C0312A0024B83F07F3991E9F21DFFFA0A3C0202B8776AC7A7C9CBFF",
INIT_13 => X"88F4C1C64044A264601144C5F1787E1C812A510885C56620590350ACD3A7D5B7",
INIT_14 => X"9054204DF56A974F92C3E20F24301300082C38C4184F10281204888298284616",
INIT_15 => X"A238CE238C8238CE238CA238CC11C6411C670C10EB4124C2B3923BF5C9710C59",
INIT_16 => X"276A11A03444922898494C5504008401230E71B3100C1634E3138C8238CC238C",
INIT_17 => X"5094650142511405194450942511425114450944519425114250144519405194",
INIT_18 => X"0944509465114251146501465014051944509445094051942501465014051940",
INIT_19 => X"2124B2DA6924965B4D5094450940519425014650142511425014450944519405",
INIT_1A => X"7DF7DF6FEFFCFDFD796ED1DCF3CF3DF6CE7F7B9DB7FF3A7E1FBC6DB7E8418A88",
INIT_1B => X"EEF77BBDDEEF77BBDDF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF",
INIT_1C => X"024F77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDD",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE056",
INIT_1E => X"5574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF80000000000000000000",
INIT_1F => X"D16AABAF7AAA8BFFAA802ABFF087FFDF5508003FEBA087FD54BA080415400555",
INIT_20 => X"AFFD54AAF7D168B45AAAABDF55AA802AA1000003FEBA00002AABA5D2EBFEBAAA",
INIT_21 => X"00003DE005555575EFA2D142145A2FFE8B45FF80001555D2E955FFFFD5421EFA",
INIT_22 => X"F5D7FC00BA5D5568AAAF7AAAAAAAAA802AABA082E954005500021FF5D2EBFF55",
INIT_23 => X"BAFFD5420AAAA843DFFFAAD1554005D7FD74AAAA840014500517FFEF007BEABF",
INIT_24 => X"4BAA2AABDE0055517FF555504154BAA2FBEAA105D2E97410FFD16AAAA5D2ABDE",
INIT_25 => X"0000000000000000000000000000000000000000000028BFF085555545550017",
INIT_26 => X"D24821E84124285C51574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7800",
INIT_27 => X"428A925D2AB8EBABEDB6AA92F7AAA8BC7B68A28BC70075FDF45080A3AEAA007B",
INIT_28 => X"2A925FFFFD1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0A38EBA1C0",
INIT_29 => X"100021FF492AB8F7D1C0438E38145B575EFA2DB45145B6F5EFB6DF78E0514555",
INIT_2A => X"55517DFC70875EABC7557FC20AA415F68AAAF7AAAAA82BE8A28A921424974004",
INIT_2B => X"0FFDB6FABA542ABAE2AF7DF470AABE8A3AFD7A2DF55400557FD54AABE84001C5",
INIT_2C => X"EF005557545490012482B6A0BAE2849043AFED1C0E10492B6FFEFA105D2A9541",
INIT_2D => X"E005D2AAABEFFB8000000000000000000000000000000000000000000000428B",
INIT_2E => X"FF55082EA8AAA087FC20105504000AA5955554BAFFAEBDE10F7FBFDEBA007BFD",
INIT_2F => X"28A00512AA8AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3AAAAB4500557",
INIT_30 => X"57FFEFFFAA97545552A821EFFBD557555AAFBC2000A2D57FFFFF7AEBFF55FF80",
INIT_31 => X"AAAAA005D04174100800021FF002EA8BEF5D0428ABA597FD55FFA2FFD5555FFD",
INIT_32 => X"D7BD54AAF7800015551517DF45005168B55557FC0012087FEAABAF7AAAAA10F3",
INIT_33 => X"FFFFFFE005D2A95410F7FFFFEBA5D2EA8ABAFBFFD74BAF7AAA8B45AAFBD54005",
INIT_34 => X"000000000000002ABEF005555555000402000FF802AAAA04452ABFF592E80010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000006000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C030028180004003220200403302301C0381A0082",
INIT_01 => X"A74041C838394848188160000C42426041000000090800090210000008510200",
INIT_02 => X"080108200C1000004465580000C0080100000000010432400800800009882050",
INIT_03 => X"080200010C234040842248600210812183806584488000103080014E88C10000",
INIT_04 => X"0040584288A6C210003120000000001002A0E8A910A072101000400A00203040",
INIT_05 => X"04096A019400C118414A00014000002014100128005004020010A0C044C02800",
INIT_06 => X"20200A301223FC029931E9931900002224240249A6D3E808D51FE00909108222",
INIT_07 => X"0008040000220001820000010C0810211A440014A040200E8240089000080002",
INIT_08 => X"0040081A08944010007FA038020080880B0104182000000000090F8102041320",
INIT_09 => X"17E2FD200240B4A409223F020888100808200450001A401BF82C21185C81744A",
INIT_0A => X"0602A0244285180542402180D001BE1907939120000020044184890800011000",
INIT_0B => X"0F0400091081190E4490A502D2A36951B428DB14A688051A5E21214601A01A22",
INIT_0C => X"455D0018101480000000A01034101480000000A01033A0081300000000001880",
INIT_0D => X"0001A0F4101480000000A01034101480000000A0103142000040000000000000",
INIT_0E => X"00000000000041E8002900018040000000000000466800C20004090000000000",
INIT_0F => X"0000034D242C2000502000000080028000000000000000240946800142000040",
INIT_10 => X"20900000001A60F0000200000000002007F000322010480000000D1A00040440",
INIT_11 => X"2018000000000025D00008958010440000000000403F4000808800000068D240",
INIT_12 => X"101280008200800000000000086670000CC0000100000000000087C000301400",
INIT_13 => X"C8B5800720849A72700094A2202301F05103202420000810C219500150002800",
INIT_14 => X"81088A454110030212C140813204D0A0888C000118471DE126805432A62A1586",
INIT_15 => X"4096C4096C2096C2096C6096C444B6004B600C446B0104D09190013589701C11",
INIT_16 => X"108D19D1804A8000904C421852240821978221B0044245B25B456C0096C0096C",
INIT_17 => X"69DA368DA1695A568DA3685A1695A768DA3685A569DA768DA1685A569DA76C5A",
INIT_18 => X"85A569DA1685A369DA5695A368DA169DA7695A168DA3695A5695A368DA3695A5",
INIT_19 => X"7638C31C71C718638E685A569DA7685A368DA5695A768DA1685A7695A168DA36",
INIT_1A => X"1C71C73B676CEDED7DE2F4DDF7DF7DF7CE7F8FF0F4FA957FCF9F7CF7F40A0010",
INIT_1B => X"FE7F3F9FCFE7F3F9FC71C71C71C71C71C71C71C71C71C71C71C71C71C71C71C7",
INIT_1C => X"2BE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"0000000000000000000000000607C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF019",
INIT_1E => X"43DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFF80000000000000000000",
INIT_1F => X"D17DEBA0855421455555574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF8",
INIT_20 => X"87FFDF5508003FEBA087FD54BA000415400550428AAAAA84021FF007BD54BAAA",
INIT_21 => X"F7AAA8BFFAAD1554BA002A95555A28417400AAFBE8ABAF7FFD54AAAA802ABFF0",
INIT_22 => X"0FFFBD5545080417555A2D17FE1000003FEBA00002AABA5D2EBFEBAAAD16AABA",
INIT_23 => X"FFFFD5421EFAAFFD54AAF7D168B45AAAABDF55AA802AA100000001EF087FEAA0",
INIT_24 => X"B45FF80001555D2E955FFFF843DEAAA2803DFEF0855401FF082EA8B555D7FC21",
INIT_25 => X"00000000000000000000000000000000000000000055575EFA2D142145A2FFE8",
INIT_26 => X"6FA92552AB8FEFF78E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FF800",
INIT_27 => X"E001EF147BD2482BED57AE921451421555551574BAB68A2DA00FFFFFFE38085F",
INIT_28 => X"FFD24BAB68A28BC70075FDF45080A3AEAA007BD24821C04124281C0E2DA82BE8",
INIT_29 => X"D2AB8EBABEDB6AA92F7AAA8BC7B6D5524AA14209557DA28E15400BEF1EFA92FF",
INIT_2A => X"5D0E071FF0071EDA38F7F1D5555000417545B6D178E281C0A38EBA1C0428A925",
INIT_2B => X"70824A8B555C7FC2147F7D1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA10",
INIT_2C => X"EFA2DB45145B6F5EFB6DF78E05145552A925FFFF8E3DE82BE8E38FFF0851401C",
INIT_2D => X"000557FE8A00F38000000000000000000000000000000000000000000005B575",
INIT_2E => X"DE10F7FBFDEBA007BFDE005D2AAABEFFBAABDFEFAAFBC00BA007BC0000FFD542",
INIT_2F => X"000AA592ABFE00F7AA821FF557FC0010F7D168A105D55421455155554BAFFAEB",
INIT_30 => X"E95410F7D57DE00FFFBC00AAFBAAAAB4500557FF55082EA8AAA087FC20105504",
INIT_31 => X"2AA8AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3D5400BA5504155EFAAA",
INIT_32 => X"7AEBFF55FF8028A00512E975FF08557FEAAF7D157545080417545F7D56AAAA59",
INIT_33 => X"F7AAAABEF005542155000028B555D7FC2145F3D557555AAFBC2000A2D57FFFFF",
INIT_34 => X"0000000000007FD55FFA2FFD5555FFD57FFEFFFAA97545552A821EFFBAABDE00",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000004800000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992006",
INIT_01 => X"A34009C0383848481C00E0000E01426040000000080000080200010000510204",
INIT_02 => X"4801082048100000446558000080000041000000000622400800000009000010",
INIT_03 => X"080001038CA14840842248400210812102000400088000003080014688800000",
INIT_04 => X"000040048106000040120000000000100220C8A5108032140004500800603000",
INIT_05 => X"04096A009000410041480081000000201000012800400022801080C0C0C82000",
INIT_06 => X"232086381A8001220021E0021803002224240248040360889100100909000222",
INIT_07 => X"0008055000220409020000090C0810211A04001420602000D2500810000C4903",
INIT_08 => X"8040491A809041100001400042409098090006102000000000010F8102041320",
INIT_09 => X"340C013102002420012200820D89140800004010900A4010002C8118D0024412",
INIT_0A => X"A221A5000800914000400888C00100200B0310200008B2066313894800631400",
INIT_0B => X"0010000800010004088105020100008000400120800000200404002450004000",
INIT_0C => X"4409081C1000000000F001F02C1000000000F001F021141A12000000000010B0",
INIT_0D => X"383480CC1000000000F001F02C1000000000F001F023420000000004C3201C51",
INIT_0E => X"00019860078641084039000000000002C0E00E0E404900E200000000000B0380",
INIT_0F => X"120C8908146000105120000000000004004160C0301D07001D04820342000000",
INIT_10 => X"000021908C4842FC000000030F000FE00600103BA0000010C8462414E8000006",
INIT_11 => X"000004C3201C60A400100DD5800000013098038D40309D000000C2419120A740",
INIT_12 => X"901A800030040902C0807C0E00C440100DDD000000411C81078884004035DC00",
INIT_13 => X"140A000410401400201020820022000250400040002211148019064200402A32",
INIT_14 => X"01889A4543148282A01415B04009904A80890033679459A926801054001C0050",
INIT_15 => X"159201592055920559205592070C901AC901A100804000801210541403C05130",
INIT_16 => X"2460010004428008904C085D44200D8001112804CDE1C483480D201592015920",
INIT_17 => X"0080200806008020000000004000020080200802000000000000000008020480",
INIT_18 => X"1000008020080000000000020080200000000000080600802008000000400000",
INIT_19 => X"5841040002082080000180200000000020180200800000000100200802000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000005428A94",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"E480000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE031",
INIT_1E => X"BC00AAF7D5575455D557DFEF002AAAB55002E820AAAA80000000000000000000",
INIT_1F => X"AEAAB55007FD74AAAA843DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFF",
INIT_20 => X"2802AA10FFFFFDE0008556AABA5D2ABFFEFFFAAAAAAAF7D57FFEFF7D555555A2",
INIT_21 => X"085542145552ABDFEFFFAA801EFFFFBFDF550000175555504175450055574AAA",
INIT_22 => X"0082A975EF00003DF55555168A00000428AAAAA84021FF007BD54BAAAD17DEBA",
INIT_23 => X"AAFF802ABFF087FFDF5508003FEBA087FD54BA000415400557BD74BAFFD14000",
INIT_24 => X"400AAFBE8ABAF7FFD54AAAAAEA8ABA55557FEAAA2843FF55A2AEA8B55AAAABDE",
INIT_25 => X"00000000000000000000000000000000000000000051554BA002A95555A28417",
INIT_26 => X"C20825D7FE8A92FFFFC70BAE3D155555415178FD7082EAAB550820870BAAA800",
INIT_27 => X"578FFFEBD55557DBEA4AFB550871D7482AA8E3DFFFAAFFD04AA415B52492B6F5",
INIT_28 => X"0E175550051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7A0ADABAEBD",
INIT_29 => X"47BD2482BED57AE921451421555524BDFD7FFA4801D7F7F5FDF55000E1754541",
INIT_2A => X"1C7BD2482E3D1450381C20905EF08003AF55415F6DA38080E2DA82BE8E001EF1",
INIT_2B => X"5BEAAAFB55ABA0BDE02EB8A28BC70075FDF45080A3AEAA007BD24821C0412428",
INIT_2C => X"AA14209557DA28E15400BEF1EFA92FFFFD24BAB6A4A8A82495F78E92AA843DF4",
INIT_2D => X"B450800174BAA680000000000000000000000000000000000000000000055524",
INIT_2E => X"00BA007BC0000FFD542000557FE8A00F3FFD54BAAAD15754508556AB45002AA8",
INIT_2F => X"AABEFFB803DEAAAAD56ABEFAAD5575EFF7803DF45085557410AEAABDFEFAAFBC",
INIT_30 => X"57FF55082E97555002E955550C55554BAFFAEBDE10F7FBFDEBA007BFDE005D2A",
INIT_31 => X"2ABFE00F7AA821FF557FC0010F7D168A105D554214551003FF45FF8400145FFD",
INIT_32 => X"87FC20105504000AA597FC2010A2D1554AA5500021EF000028B55087BFDEBA04",
INIT_33 => X"007FE8A00A2803FF45F7AABDF55AA843FE10AEAAAAB4500557FF55082EA8AAA0",
INIT_34 => X"00000000000055400BA5504155EFAAAE95410F7D57DE00FFFBC00AAFB8028A00",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"A140084000080048040100000202026040000000180800080200010048510204",
INIT_02 => X"080108000090000004655C000080000051000000000402400800000009000010",
INIT_03 => X"0000000100300C40842240000210810002800584488000103080894288800000",
INIT_04 => X"0002584280A2C21000110300100000100220C8C910A032541000090A00643000",
INIT_05 => X"04092A001400D100410A002140004020140001A9005000004810A1C0044D2800",
INIT_06 => X"0360000010EFFD229911C9911820002080258A09A2D3E102137FE0094910A222",
INIT_07 => X"0000004000220400120000090C0810210A040034A040000046180810000C4907",
INIT_08 => X"80404050D88C24510001400042008088090004012000000000010F8102041320",
INIT_09 => X"20080120024030A4090200828C880208002044C0843B44100228A1585C81740A",
INIT_0A => X"142180860A84802042C82180D0010039039390200008B20E2300086800400640",
INIT_0B => X"003000091084190644810502D0A16850B4285B14A688011A1409212008F05E20",
INIT_0C => X"400104080010001E0FF00010000010001E0FF0001002200A1300000000000080",
INIT_0D => X"000080000010001E0FF00010000010001E0FF000100440000040F517CF600000",
INIT_0E => X"E587F9E000004008100800008000ED0FC7E000004000804000000809963F1F80",
INIT_0F => X"36000100202C0020100000000802419660CFE7C0F00000000800810040000040",
INIT_10 => X"0618E7B0000800000003F80FFF0000200018021000030C73D80004000000585F",
INIT_11 => X"078A8FCF600000201802008001006AA3F1F80000400000000B0BD6C000200000",
INIT_12 => X"0041120370DCAD1FC18000000040180200800005D5C3FD800000806008100000",
INIT_13 => X"48A480072284983230101402200200111103202420000880C218000150100800",
INIT_14 => X"2B888A4500048240C08400843204502000890001000415E12480003002944281",
INIT_15 => X"0480004800048000480004800004002240020854884000901212140011C01079",
INIT_16 => X"346D19D1A4C08028904C4E1D7224086590800420044040020004004480004800",
INIT_17 => X"68DA368DA368DA368DA368DA368DA1685A1685A1685A1685A1685A168DA36CDA",
INIT_18 => X"8DA3685A1685A1685A1685A368DA368DA368DA3685A1685A1685A1685A1685A1",
INIT_19 => X"40000000000000000068DA368DA368DA1685A1685A1685A1685A368DA368DA36",
INIT_1A => X"3CF3CF6FE23CCD8D00A281F5B2DB2CA78A543EBC57A10A245DA975D640088884",
INIT_1B => X"3E1F0F87C3E1F0F87CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"5DA9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0F87C",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00B",
INIT_1E => X"40000000043DF55087BC01EF007FD75FFFF84000AAFF80000000000000000000",
INIT_1F => X"2EBFE10A28028AAAAAFBC00AAF7D5575455D557DFEF002AAAB55002E820AAAA8",
INIT_20 => X"2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFAA95545552ABFE00087BC00AA08",
INIT_21 => X"007FD74AAAAD57FF45002A975FF007BE8BFFA2FBFFFFFAAD5400AAFF843DFEFA",
INIT_22 => X"5AAFBE8A00082A97410F7D5555EFAAAAAAAAAF7D57FFEFF7D555555A2AEAAB55",
INIT_23 => X"450055574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFFAA8200055555554",
INIT_24 => X"F55000017555550417545000015545087BC2010AAD54014500516ABFFA2AABDF",
INIT_25 => X"0000000000000000000000000000000000000000002ABDFEFFFAA801EFFFFBFD",
INIT_26 => X"AAB550820870BAAA8407000140038F450075C71FF087BD75D7FF84050BAEB800",
INIT_27 => X"AB8E10007FC50BA002ABFE00AA8A2AABABEFFC70BAE3D155555415178FD7082E",
INIT_28 => X"DB45082EB8E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFA497545552",
INIT_29 => X"BD55557DBEA4AFB550871D7482AAD17DF451C24955EF0875EFBD7B6F1FFFC7BE",
INIT_2A => X"F7AA87000415B5057DAAFBE8A10082092410EBD5505EFB6A0ADABAEBD578FFFE",
INIT_2B => X"D005B6ABC7B6AABFFED0051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEF",
INIT_2C => X"D7FFA4801D7F7F5FDF55000E17545410E17555000E17545007BC0000BED14217",
INIT_2D => X"555F784174AAA280000000000000000000000000000000000000000000024BDF",
INIT_2E => X"754508556AB45002AA8B450800174BAA684174105D042AB550055555FF007BD7",
INIT_2F => X"E8A00F384175555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7FFD54BAAAD15",
INIT_30 => X"57DF55FFD57DF55FFFBD5400A2AABDFEFAAFBC00BA007BC0000FFD542000557F",
INIT_31 => X"803DEAAAAD56ABEFAAD5575EFF7803DF45085557410AED17FF455D04155FF005",
INIT_32 => X"07BFDE005D2AAABEFFBAE97410087BC21EFA2FFEAA00000002010A2D5421FFFF",
INIT_33 => X"087BC0010FFD1401EF087FE8B55FFAEBDFEF0855554BAFFAEBDE10F7FBFDEBA0",
INIT_34 => X"000000000000003FF45FF8400145FFD57FF55082E97555002E955550C2E95555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000002000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000006",
INIT_01 => X"0000098218302849180060000C004260413C0A61590001D90213C80000110200",
INIT_02 => X"680108220010000054400C00008000004100000001200240080080000908A011",
INIT_03 => X"000A0000040020400002021000000008428065044880001030818C0008C10000",
INIT_04 => X"00005042882A8210003000000800001000806080100040140080040800003140",
INIT_05 => X"0400000840000098410800010001002000000000004000002010000040002000",
INIT_06 => X"03600810100001220911E0911902000020200200A253E8000C0010080800004C",
INIT_07 => X"000408C0002204400200000B080000010C040004A0400000C0000810000C5901",
INIT_08 => X"000008002A84300000014000C2008088090008002000000000030F8000001220",
INIT_09 => X"0008012100000200001200820888010800200000000840100028800004801440",
INIT_0A => X"000090220000040400480000D0010009049090200008B2022384800802010000",
INIT_0B => X"001000090001090A4C81240050A328519428CA14328C840A5820000101500400",
INIT_0C => X"00510008100400000000A00000100400000000A00000000A12000000000000B0",
INIT_0D => X"00012000100080000000A00000100080000000A0000540000000000000000000",
INIT_0E => X"00000000000000A8000900010000000000000000060000420004000000000000",
INIT_0F => X"0000024000240000102000000080000000000000000000240000800140000000",
INIT_10 => X"0080000000120CFC000000000000000001280013E010000000000900F8040000",
INIT_11 => X"2000000000000001480006D5801000000000000000091F0000800000004807C0",
INIT_12 => X"901A800080000000000000000820080006DD000000000000000002A00019DC00",
INIT_13 => X"0200800522C01252501086222082000010012024200000048019502000000C32",
INIT_14 => X"0080004501000200089400005200D0820008000000104C4800010600BC228404",
INIT_15 => X"0001040010000104001000010440080000822900000000801010500A13404111",
INIT_16 => X"32851951A0CA8080924C06403600086491900224002200400440104001040010",
INIT_17 => X"284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A128CA328CA",
INIT_18 => X"84A1284A1284A1284A1284A328CA328CA328CA328CA328CA328CA328CA328CA3",
INIT_19 => X"10000000000000000028CA328CA328CA328CA328CA328CA328CA1284A1284A12",
INIT_1A => X"69A69A250B61004055CD1439248209070CCCF48DE68A8900401038E2550A0010",
INIT_1B => X"341A0D068341A0D068A28A28A28A28A28A28A28A28A28A28A28A28A29A69A69A",
INIT_1C => X"56C1A0D269341A0D068349A4D068349A4D068341A0D269341A0D269341A0D068",
INIT_1D => X"0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE052",
INIT_1E => X"57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D00000000000000000000",
INIT_1F => X"D1575EF00557DF555D040000000043DF55087BC01EF007FD75FFFF84000AAFFD",
INIT_20 => X"7D5575455D557DFEF002AAAB55002E820AAAA843DFEF00517DEBA007BFDFEFFF",
INIT_21 => X"A28028AAAAAAABDF45F7803FFEF555568AAAF7802AA00FFFBD7555087BC00AAF",
INIT_22 => X"5087BD54BA550417400085155555082A95545552ABFE00087BC00AA082EBFE10",
INIT_23 => X"555D043DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00AA552E9554",
INIT_24 => X"BFFA2FBFFFFFAAD5400AAFF8402000A2FFFDF555D7BE8BFF5D51575EFA280175",
INIT_25 => X"000000000000000000000000000000000000000000557FF45002A975FF007BE8",
INIT_26 => X"D75D7FF84050BAEBDF78F45B68010482415B471C7E3DF451EFBEFBFAF4549000",
INIT_27 => X"17DE82007FFAFEFE3DB505EF1C5B7AF45490407000140038F450075C71FF087B",
INIT_28 => X"FFD55451C7FC70BAE3D155555415178FD7082EAAB550820870BAAA8438FFF005",
INIT_29 => X"07FC50BA002ABFE00AA8A2AABABEAEB8F45F78A3DFD741516DAAAE38E2DA28EB",
INIT_2A => X"FFFFC20BA5D2E905550071D54825D0A1543808515756D1C2497545552AB8E100",
INIT_2B => X"F5D55505FFBE801256D490E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92",
INIT_2C => X"451C24955EF0875EFBD7B6F1FFFC7BEDB45082EB8002000AAFFFDF6D417FEABE",
INIT_2D => X"5EFF7FBE8B5500000000000000000000000000000000000000000000000517DF",
INIT_2E => X"AB550055555FF007BD7555F784174AAA2FBEAB45F78402010007BD5545AAFFD5",
INIT_2F => X"174BAA68028BEF00517FE10007BE8BFFAAFFC01FF557FE8B550004174105D042",
INIT_30 => X"57FEAAAAAEBFEAAAAFFD5545557FD54BAAAD15754508556AB45002AA8B450800",
INIT_31 => X"04175555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7AAAAB45F7AEBFF45085",
INIT_32 => X"FD542000557FE8A00F3FFC00BA552E80145005557400552A954BA0051575EF55",
INIT_33 => X"A2FBFDFFF007FE8BFF5551401EFF784021FF002ABDFEFAAFBC00BA007BC0000F",
INIT_34 => X"000000000000517FF455D04155FF00557DF55FFD57DF55FFFBD5400A28400010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000004000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A14009801830084C182060000C10424840000000080000080200000000110204",
INIT_02 => X"0801080200100000046558040080000041000000002402400800000009008010",
INIT_03 => X"00020201040000D0842242024210810802006400088000003080054288C10000",
INIT_04 => X"0000400088020000003020002000001002A0E881108032100002000800203040",
INIT_05 => X"04092A081000411841480001000000201000012800400010001081C040402000",
INIT_06 => X"03600810100001220001E0001802002020240208000369001500100909000266",
INIT_07 => X"0000004000220440020000090C0810210A040004A0410000C0000810000C4901",
INIT_08 => X"0040480000802100100140004200808809000C002000000000010F8102041320",
INIT_09 => X"2008012000000000000200828888800808000410800840100220211850004442",
INIT_0A => X"040180240A80800442400004C0010000060210200008B2022304880800010000",
INIT_0B => X"0030000000010008008020020100008000400120800004004821202001A05A00",
INIT_0C => X"40510008101480000000A01004101480000000A0100000001300410402080080",
INIT_0D => X"0001A004101480000000A01004101480000000A0100540000040000000000000",
INIT_0E => X"00000000000040A8000900018040000000000000460800420004090000000000",
INIT_0F => X"0000034000082000102000000080028000000000000000240800800140000040",
INIT_10 => X"20900000001A00000002000000000020013000100010480000000D0000040440",
INIT_11 => X"2018000000000021500000800010440000000000400900008088000000680000",
INIT_12 => X"000000008200800000000000086010000080000100000000000082C000100000",
INIT_13 => X"000080000004924040008020000200101100004000000000C019500050000800",
INIT_14 => X"2B088A4541008240001000804000108280800001001051A12481041080801010",
INIT_15 => X"4480004800048004480044800044000240022100884000901210440003C14110",
INIT_16 => X"06E00000044200009849485D4020080000140004046240020044000480044800",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802000000400",
INIT_18 => X"0000000000000000000000020080200802008020080200802008020080200802",
INIT_19 => X"1000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"1451451AA654199951A24454514514F0CA940FE0D39712615FAD555204428290",
INIT_1B => X"CA6532994CA65329945145145145145145145145145145145145145145145145",
INIT_1C => X"670E572994CA6532994CAE572B95CA6532994CA6532B95CAE572994CA6532994",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE01C",
INIT_1E => X"03FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF0800000000000000000000",
INIT_1F => X"7FFDF45FFFBC2010AAD57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D0",
INIT_20 => X"0043DF55087BC01EF007FD75FFFF84000AAFF8002155AAFFE8B45AAD54000008",
INIT_21 => X"00557DF555D517FEBA082A801EFF7FBD5400FFD568B555D00155EF0804000000",
INIT_22 => X"AF7FBFDE00A2FBC0145005168A10AA843DFEF00517DEBA007BFDFEFFFD1575EF",
INIT_23 => X"EF5D7BC00AAF7D5575455D557DFEF002AAAB55002E820AAAA803FEBA082AAAAA",
INIT_24 => X"AAAF7802AA00FFFBD7555082E82155FFAEAAB55AAD568B455D00154BAFFFBD75",
INIT_25 => X"0000000000000000000000000000000000000000002ABDF45F7803FFEF555568",
INIT_26 => X"451EFBEFBFAF4549003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC700000",
INIT_27 => X"5EDB6DAADF470280075FFF45E3F1C7038A2DF78F45B68010482415B471C7E3DF",
INIT_28 => X"0A175C7000407000140038F450075C71FF087BD75D7FF84050BAEB8002155BEF",
INIT_29 => X"07FFAFEFE3DB505EF1C5B7AF45495B7DEAA0824851EFEBFBD2410EBD168B7D41",
INIT_2A => X"AA8038EAA0824A8AAAEBF5FAE28AAF1C2155005F68A10A28438FFF00517DE820",
INIT_2B => X"D4104104AAF7F1D75EF557FC70BAE3D155555415178FD7082EAAB550820870BA",
INIT_2C => X"45F78A3DFD741516DAAAE38E2DA28EBFFD55451C2087155EBA4A8B7DAADF68B7",
INIT_2D => X"FEFA2AEAAB55000000000000000000000000000000000000000000000002EB8F",
INIT_2E => X"2010007BD5545AAFFD55EFF7FBE8B5500043FE00F7D17FEBAA2D5574BAAAD17D",
INIT_2F => X"174AAA28002155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAB45F7840",
INIT_30 => X"BC2000AAD16ABFF002A975450004174105D042AB550055555FF007BD7555F784",
INIT_31 => X"8028BEF00517FE10007BE8BFFAAFFC01FF557FE8B55007FFDEAA0004175FFA2F",
INIT_32 => X"02AA8B450800174BAA68428AAA08042AABAAAD56AABAAAD140155087FEAA10A2",
INIT_33 => X"A2842ABEFAAFBE8BFF0004020AAFFD5555EF557FD54BAAAD15754508556AB450",
INIT_34 => X"0000000000002AAAB45F7AEBFF4508557FEAAAAAEBFEAAAAFFD5545550015555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000047FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B83008481800E0000C26426040000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"00080D4912E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"000048048002400048150000000002504230C899109032100020160880223000",
INIT_05 => X"040B2A229100410041088011100022201200012840440000B01088C0005C2400",
INIT_06 => X"03286A287E4003225021C5021880C02000A40249048363A5990010090908022A",
INIT_07 => X"8320694044222987020C80152D8910210A0400252B74200045C86810000C5B05",
INIT_08 => X"00404126509804400501400242C0B0B83B0134702000000000191FA162841324",
INIT_09 => X"2008013002000220001240820F8B2A08000040409018401001200159D80D64AA",
INIT_0A => X"91019B02080885200042E098C00101B0070310200008B60A23A51B2802067327",
INIT_0B => X"003000080802500C088325828102408120409120940680100504022148504440",
INIT_0C => X"1501D5761B011986695014A96E1A8119865A5018C5A0A00012004104020808B0",
INIT_0D => X"A2600AAE1A811986695014A96E1B0119865A5018C5AF0062C38A4DB680A0D824",
INIT_0E => X"1DB528802CAB184E8F4101621B1BAC845542056A289A1BB2078A922DA2A8B180",
INIT_0F => X"7A3D94392000224ACDE215883078681B5C05AA429189B60AC43CEC7F0272C384",
INIT_10 => X"134CD551BCA1C90006C0C2958502861120C003104289A668B8CAB27010633831",
INIT_11 => X"82806CA64090B89E015AAA880E48382EB8804B020A06020C67061BC785938085",
INIT_12 => X"470126C6284B2D20410AB4503089C00A8280819A5539D503336D61056ABA0062",
INIT_13 => X"000080060040142020015001004A00080042004000E8089C9003066E03513E41",
INIT_14 => X"010CBA45367082014000908020349320008000A1000C09A9348498B000000000",
INIT_15 => X"C32A0832A0C32A0C32A0832A0C19504195040040000000801010028001400010",
INIT_16 => X"2468118104400000904C0C0964200841010954000444D280140050C32A0832A0",
INIT_17 => X"4090240902409024090240902409024090240902409024090240902409024090",
INIT_18 => X"0100401004010040100401024090240902409024090240902409024090240902",
INIT_19 => X"0000000000000000004010040100401004010040100401004010040100401004",
INIT_1A => X"410410502A441495418984700000005088804180C0B10A04D0A7104201400284",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000010410410",
INIT_1C => X"7800000000000000201000000000000000000008040000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE060",
INIT_1E => X"4155EFAA842ABEFA280155EFFFFBC01EF0855400005500000000000000000000",
INIT_1F => X"FBFFF4508514000000003FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF080",
INIT_20 => X"280154BA5555401EFFFD5421EFA2FFFFF555D51575FFA2FFD75FF550015400FF",
INIT_21 => X"FFFBC2010AAD568AAAAAD142145FF80155EF0051555FF0804155FFF7D57DF45A",
INIT_22 => X"008001540008514215555003DFFFA28002155AAFFE8B45AAD540000087FFDF45",
INIT_23 => X"0000040000000043DF55087BC01EF007FD75FFFF84000AAFF802ABFFA2AABFE1",
INIT_24 => X"400FFD568B555D00155EF085168B45085142010FFAE800AA5D7BFDF45F7FFEAA",
INIT_25 => X"000000000000000000000000000000000000000000517FEBA082A801EFF7FBD5",
INIT_26 => X"7DF7DA2AEB8FC70000175EFB6802DBC7BE8A155EFE3FBC71FF145B4203855000",
INIT_27 => X"5D05EF550E15400E3F1FFF7D085B420381C003DE10BEF5EDAAAAAD547038EBD5",
INIT_28 => X"04105C7F7DF78F45B68010482415B471C7E3DF451EFBEFBFAF45495F575FFBEF",
INIT_29 => X"ADF470280075FFF45E3F1C7038A2DB68ABAB6D145145FF84155D7085B555C714",
INIT_2A => X"EB8428BEFBEA4BDE28140A1543800514515549003FFC7BE8002155BEF5EDB6DA",
INIT_2B => X"2417FFFF7DE3F1EFA10140407000140038F450075C71FF087BD75D7FF84050BA",
INIT_2C => X"AA0824851EFEBFBD2410EBD168B7D410A175C7005B6DB55145140000FFAE8508",
INIT_2D => X"5EF557BC20AA5D0000000000000000000000000000000000000000000005B7DE",
INIT_2E => X"FEBAA2D5574BAAAD17DFEFA2AEAAB550004175FFF7803DF45FFAE955EFAAFBD5",
INIT_2F => X"E8B55007FD75FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D043FE00F7D17",
INIT_30 => X"015555007FD5545550400145FFFBEAB45F78402010007BD5545AAFFD55EFF7FB",
INIT_31 => X"8002155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAAAAFFD555545FF8",
INIT_32 => X"07BD7555F784174AAA2842ABEFFF803DEAA5D2E974AA00515754500003FF55FF",
INIT_33 => X"555540000FFAE97410007BFFFFFA2D57FE105D04174105D042AB550055555FF0",
INIT_34 => X"0000000000007FFDEAA0004175FFA2FBC2000AAD16ABFF002A97545007FFFF45",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000004000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C048000C048400380000007024040000000080000088200002802153231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"421A0A0012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"02004000890200001837800001998C31C090609C104000102002140900003548",
INIT_05 => X"0402002BC200009841090001200006200800000020480010A4100100001C2000",
INIT_06 => X"033432287FC003230001D0001806C0060CB0622000037085C800100C0C200008",
INIT_07 => X"135038CE64B663DFA314C803292140890C0601F472D1640051F80C10020C493F",
INIT_08 => X"00000167C081000011814004C20481A92940EA7A3020480000071F846890162E",
INIT_09 => X"D40C01240008000080024082488BAF08000020000208401004300421800F04F8",
INIT_0A => X"F9F80FA0200E0BF40063FF9DC0010000180018200408B27E234913E900067F04",
INIT_0B => X"001100002002801000A04200000000000000000000029D204B7C0382FD0100F3",
INIT_0C => X"9628F97E0B348EDAC3900F6EFA0B158EDA93900F6EE230381208008001007A80",
INIT_0D => X"EAE64BCA0B158EDAC3900F6EFA0B348EDA93900F6EE8421392C96B1237E0D8BD",
INIT_0E => X"4CAEAD412EDD2B47CFF812A383430C669E622DBC31D73F6006A5891533EF9500",
INIT_0F => X"2E19B8BA30E022DAD8C100CA39E8CEBE66C2B083798D341B10DE7E14400392C7",
INIT_10 => X"32966471A9C5DD00B12728D5360234D62A49FAB442994B3238D4E2FB10463665",
INIT_11 => X"F0FABAC800DA550C29F36A8A2554E48A6430469392526208C6CC95C33717D885",
INIT_12 => X"2B416A51B60585A5C28895962502E9F36A828C4999AF580395542D27CDBA0020",
INIT_13 => X"0000800000001E404011F066000A000EE040000000873FB80B8A00EF03F56CC1",
INIT_14 => X"2284304D667C06CC6816B300403C13E2000000460010400000010CE080801010",
INIT_15 => X"872F0872F0C72F0872F0872F0C597863978421000800209010104ACA03414110",
INIT_16 => X"01000000104280009048004000000800001D5E05182493C5BC5AF0872F0C72F0",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0802008020080200802008000000000000000000000000000000000000000000",
INIT_19 => X"1000000000000000000080200802008020080200802008020080200802008020",
INIT_1A => X"492492240F010000146E502D4514510246088881360A95118B120CB054420210",
INIT_1B => X"6432190C86432190C82082082082082082082082082082082082082092492492",
INIT_1C => X"7FEB2592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2590C8",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"5421FF00042ABEFFF8400010082EAABFF55002ABEF0800000000000000000000",
INIT_1F => X"002ABEFFFFBD54000004155EFAA842ABEFA280155EFFFFBC01EF085540000555",
INIT_20 => X"AFBE8AAAA2D540000F7D57DF55A2AABFFEF08556AA10000028AAAFFD15541000",
INIT_21 => X"085140000005168AAA087BFFFFF5D04001FF00041554555557FE005D003FE10A",
INIT_22 => X"F0851555FF082AA8B55F7AEA8BEF5551575FFA2FFD75FF550015400FFFBFFF45",
INIT_23 => X"10AAD57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D0000145082E955F",
INIT_24 => X"5EF0051555FF0804155FFF7842AA100000020BAAA801541055042ABEFFFFBD54",
INIT_25 => X"0000000000000000000000000000000000000000005568AAAAAD142145FF8015",
INIT_26 => X"C71FF145B42038555F401D71C0A2DBC7EB80000280824ADBD7490E28BEF08000",
INIT_27 => X"A2DA82FFDB5243800002FBD7EBFBD24101C00175EFB6802DBC7BE8A155EFE3FB",
INIT_28 => X"5B7AE1041003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7005F6AA381C0",
INIT_29 => X"50E15400E3F1FFF7D085B420381C5B6AA82147FF8FEF410E001FF000E1755555",
INIT_2A => X"49000017D142E905EF1451525C7082AADB45F7AEA8BEF555F575FFBEF5D05EF5",
INIT_2B => X"041002FBEFEBFBD2410AADF78F45B68010482415B471C7E3DF451EFBEFBFAF45",
INIT_2C => X"BAB6D145145FF84155D7085B555C71404105C7F7842FA381C0A00082AA8A1041",
INIT_2D => X"F55002AA8BEF000000000000000000000000000000000000000000000005B68A",
INIT_2E => X"DF45FFAE955EFAAFBD55EF557BC20AA5D7BC01555D2EBFF55A284000AA08003F",
INIT_2F => X"AAB55007BE8AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D04175FFF7803",
INIT_30 => X"E821FF082A97555557FE8A0000043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AE",
INIT_31 => X"7FD75FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D7BE8A005D7FEABFF002",
INIT_32 => X"AFFD55EFF7FBE8B550004001FF5D2A801EF5D5142145082EBFF55F7AAAABEF5D",
INIT_33 => X"552A82010A2AA8000008043FFFFA2FBC2010A2FBEAB45F78402010007BD5545A",
INIT_34 => X"0000000000007BEAAAAFFD555545FF8015555007FD5545550400145FF843DEAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400986B830E84D182260000C1042684001000008220008A20019080A510200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00020201926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"00104884880A4400403003005800027102A0E8C110D83210642EA809C0203040",
INIT_05 => X"04092A08138041184109C001380000201A008128044E00754010C9C192D82400",
INIT_06 => X"032C7E201800012372A1D72A180000204024024954A3670819001009092C0222",
INIT_07 => X"0164004000220B40020C80052C0A12292A040005715540015E006810001C4B01",
INIT_08 => X"0040549032881001140140024200808839005C002010800000155F8122851320",
INIT_09 => X"6008012C80481284881280825A988008000040808629441005B3071859006442",
INIT_0A => X"0001B0200810940400720005C0030192072310200028B6022346080802E001A5",
INIT_0B => X"003000206822F20CA8826AC2A14250A128509528954404144C20042501004000",
INIT_0C => X"03D404A41AA5B7344C10B383081BA4B7341C10B3831034081200000000000430",
INIT_0D => X"5A2B2C381BA4B7344C10B383081AA5B7341C10B383110218CB0E54C2EA404A4F",
INIT_0E => X"3548B3A008E730A01AB113A5524E6ACA678001CE3E20A5B284ED1132909C7288",
INIT_0F => X"0A3C066430202021252991C22C99731014AC3CC0C0B8182597A801610218CB0C",
INIT_10 => X"A5C8825194332B018A444AEA2701288A15A151EC5952E44128CA194517354C18",
INIT_11 => X"635232D50048A411C158BB0A7910142C771804C8A0ADA2E6A983014780CA28B2",
INIT_12 => X"6E4023F8BE8E3E1E0109472C3EB50158BB02D09852745F80112C428562EE0353",
INIT_13 => X"00008002414032646000826080C20001104240480068001C9B9150A000029704",
INIT_14 => X"1118BA4510008241C80290882400908000A000A1000809A93485D61000000000",
INIT_15 => X"40000000000000040000000000000020000000040000008010122A8201410058",
INIT_16 => X"246A10A1044101A89A4D0C096420184321040002844840000000004000000000",
INIT_17 => X"5094250942509425094250942509425094250942509425094250942509425094",
INIT_18 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_19 => X"0000000000000000005094250942509425094250942509425094250942509425",
INIT_1A => X"75D75D7FEDFDFDFDFBEEF9DD555555F7EEFF3F7DF7FF3E7E1FBF7DF7E24502A8",
INIT_1B => X"FAFD7EBF5FAFD7EBF5D75D75D75D75D75D75D75D75D75D75D75D75D75D75D75D",
INIT_1C => X"7FEFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F780000000000000000000",
INIT_1F => X"AA97400AAD540155A2D5421FF00042ABEFFF8400010082EAABFF55002ABEF085",
INIT_20 => X"A842ABEFA280155EFFFFBC01EF08554000055043DEBAF7843FFFFF7AABDF55A2",
INIT_21 => X"FFFBD5400005568A1055043DEBAAAFFE8B45557FD7410552EAAABAAA84155EFA",
INIT_22 => X"AA2FFE8ABAAA8428A00087BD7555FFD56AA10000028AAAFFD15541000002ABEF",
INIT_23 => X"55A2803FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF085557545FFD17DEB",
INIT_24 => X"1FF00041554555557FE005D0000155557BEAABA5D2ABDF450851420AA5D7FD55",
INIT_25 => X"0000000000000000000000000000000000000000005168AAA087BFFFFF5D0400",
INIT_26 => X"ADBD7490E28BEF08516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EB800",
INIT_27 => X"03FFD7EBA4BDF45AAAA90410BEDF45155A2DF401D71C0A2DBC7EB80000280824",
INIT_28 => X"2AAFA82B680175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550E38E92EB8",
INIT_29 => X"FDB5243800002FBD7EBFBD24101C556FA38490A3FE92BEFFEAB45417FD24385D",
INIT_2A => X"00515056DE3D17FE92BEF1EFA92AA8428A10007FD557DFFDF6AA381C0A2DA82F",
INIT_2B => X"5085B400925D7FD557DA2803DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7",
INIT_2C => X"82147FF8FEF410E001FF000E17555555B7AE10410E00155497FEFABA4120B8F5",
INIT_2D => X"ABAA2FBD7545AA8000000000000000000000000000000000000000000005B6AA",
INIT_2E => X"FF55A284000AA08003FF55002AA8BEF00517FE00082EBDF45AA8428A10085568",
INIT_2F => X"C20AA5D2EA8A00A2803DF45AA843DF55AAAE82000F7FBD5545AAFBC01555D2EB",
INIT_30 => X"FE8B55087FC00BA552ABFE10F784175FFF7803DF45FFAE955EFAAFBD55EF557B",
INIT_31 => X"FBE8AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D517FEAA082EBFE10F7F",
INIT_32 => X"AD17DFEFA2AEAAB550051401FFA2D57FE10F7D57DE00AA842AA00007FD75FFF7",
INIT_33 => X"007BFDEAA08042AB45087FC0010557FD55FFAA843FE00F7D17FEBAA2D5574BAA",
INIT_34 => X"0000000000007BE8A005D7FEABFF002E821FF082A97555557FE8A00002E82155",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000067FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"0002074F200904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000480488024000403000000000001002A0E881108032100002000800203040",
INIT_05 => X"04092A081000411841080001000000201000012800400010001081C000402000",
INIT_06 => X"033D7880500001221021C1021800002000240249048361001100100909000222",
INIT_07 => X"9020304000220050020480152D0A142D0A8400043B45400040006810000C5901",
INIT_08 => X"0040400010880000100140024280808829029C002000000000053FA142051324",
INIT_09 => X"6008012000000000000200820888800800004000800840100020011858006442",
INIT_0A => X"000110200800840400400005C0010190070310200008B202236D080802000001",
INIT_0B => X"003000000000100C088020028102408120409120940404104C20002101004000",
INIT_0C => X"2050805210040000B0E0A0000210040000E0E0A0000190081200000000000000",
INIT_0D => X"0111300210008000B0E0A0000210008000E0E0A0000B02740421A0E5D1A02400",
INIT_0E => X"C0715C40110080A4006110510C14D18178E01200860008920106460D4501CB00",
INIT_0F => X"500002411420220080220C0093C38923240ABBC00905C33C6000400F02740412",
INIT_10 => X"9682398000120800658992F3C700C3018120000041DB011CC000090012565306",
INIT_11 => X"B7A0B1E240240A8340000200067EAA8CB65809240C09024A4AE0CA0000480083",
INIT_12 => X"00845C7DB0D0200900422ACA4B28000002002B46867DBC002A830280000800F7",
INIT_13 => X"000080020040126060008020000200000042004005800004801150A003412440",
INIT_14 => X"01088A4500008240000000802000908000800001000009A92481041000000000",
INIT_15 => X"0000000000400000000000000400000000000000000000801010000001410010",
INIT_16 => X"246810810440000090480C096420084101040000044040000000004000040000",
INIT_17 => X"4090240902409024090240902409024090240902409024090240902409024090",
INIT_18 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_19 => X"0000000000000000004090240902409024090240902409024090240902409024",
INIT_1A => X"3CF3CF3FE77DDDDD55E6D5FCF3CF3DF7CE5C8FF0F7BE9D75CF9F7DF650400280",
INIT_1B => X"FE7F3F9FCFE7F3F9FCF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"8007F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE07F",
INIT_1E => X"17DF45AAD157400007BEAAAAAAAE955555D5568A105D00000000000000000000",
INIT_1F => X"AA800AAF784020AAF7D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7D",
INIT_20 => X"0042ABEFFF8400010082EAABFF55002ABEF085155400FFD1420100055574AAA2",
INIT_21 => X"AAD540155A28028B550051574005D7FFFE105D7BD7545A284020BA0055421FF0",
INIT_22 => X"00851421FF5D7FFDEBA085168B45FF843DEBAF7843FFFFF7AABDF55A2AA97400",
INIT_23 => X"FF5504155EFAA842ABEFA280155EFFFFBC01EF08554000055002AB455D514201",
INIT_24 => X"B45557FD7410552EAAABAAA8017400AAD140000002EBFFEFA2AAA8BEFF780021",
INIT_25 => X"0000000000000000000000000000000000000000005568A1055043DEBAAAFFE8",
INIT_26 => X"F8E38E3DF45155EBD17FF6DAADB504001C71EDA82AAA0955455D556DA0049000",
INIT_27 => X"B420101C55554AAAAA480082FF84000BAEBD16DA82410A3FFD7AAA4B8E824971",
INIT_28 => X"8405092085F401D71C0A2DBC7EB80000280824ADBD7490E28BEF085157428FFD",
INIT_29 => X"BA4BDF45AAAA90410BEDF45155A28E2AB7D0051504005D71F8E004975D556DB6",
INIT_2A => X"550028B6D5D51420101C5B401EF417BFAEAA08516AB45E38E38E92EB803FFD7E",
INIT_2B => X"7A2AEAFBC7EB80071FF5500175EFB6802DBC7BE8A155EFE3FBC71FF145B42038",
INIT_2C => X"38490A3FE92BEFFEAB45417FD24385D2AAFA82B68015400AADB40000082EBFFC",
INIT_2D => X"54555557FE1000000000000000000000000000000000000000000000000556FA",
INIT_2E => X"DF45AA8428A10085568ABAA2FBD7545AAD17DFFFAAFFC200055557DE00A28015",
INIT_2F => X"A8BEF0051554AAFFFFC00105D55554BAA28400000F784020BAAAD17FE00082EB",
INIT_30 => X"568A000051575FFF78415410087BC01555D2EBFF55A284000AA08003FF55002A",
INIT_31 => X"AEA8A00A2803DF45AA843DF55AAAE82000F7FBD5545AAAEAABFF0051400105D5",
INIT_32 => X"AFBD55EF557BC20AA5D042ABFF555142000557FC01EF007FEAABA00556AB55A2",
INIT_33 => X"A2FBC0010082EBDF55A2AABDF45A284175FF5D04175FFF7803DF45FFAE955EFA",
INIT_34 => X"000000000000517FEAA082EBFE10F7FFE8B55087FC00BA552ABFE10F78415400",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000100000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"000440009282000001100000000000100220C8811080321000000228002A3000",
INIT_05 => X"04092A0010004300418800510000A6201000012A64400000145080C000422000",
INIT_06 => X"032B1800100001220001C00018821020402402080003772019001009090002AA",
INIT_07 => X"0000004000220000021840010C8912250A0400042044400040006810000C4901",
INIT_08 => X"0040400022810000058140024280A0A8190004002030C00000016F8122041320",
INIT_09 => X"E0080120000000000002C0820888008800000000800840100020011850004402",
INIT_0A => X"00013000080094000062000180010180060210200008B2022304080800000003",
INIT_0B => X"0030000000000008008020020000000000000100800000000000002500004000",
INIT_0C => X"0000000010108000000000000010108000000000000230001200000000000420",
INIT_0D => X"0000000010140000000000000010140000000000000100000040000000000000",
INIT_0E => X"0000000000000000000100008040000000000000000000020000090000000000",
INIT_0F => X"0000000030002000406000000000068409014000000000000000000100000040",
INIT_10 => X"2010000000000800000201000800000000000000400048000000000010000440",
INIT_11 => X"00184400A0000000000002000000441108800000000002008008000000000080",
INIT_12 => X"0000000242038B82800000000000000002000001000000000000000000080000",
INIT_13 => X"000080000000100000000005C04A000000400000000000000001062000000400",
INIT_14 => X"01088A4500008200000000800000100000800001000001A12480001000000000",
INIT_15 => X"4000040000000000000000000400002000020000000000801010000041400010",
INIT_16 => X"0460000004400000904808094020080000000000044040000000004000040000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000400280",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FC00000804154AA5D00001EFF78428AAA007BC2145F780000000000000000000",
INIT_1F => X"55400AA007FC2000F7D17DF45AAD157400007BEAAAAAAAE955555D5568A105D7",
INIT_20 => X"D043FFFFAAAABDEAA557BFDE00FFD140155F7FBD74AAAAD17DF45F7D1421EF00",
INIT_21 => X"F784020AAF7FFFDF45FF84000BA552ABDFEF08517DF55A2FBEAB555D556AAAA5",
INIT_22 => X"5AAFFEAB45F7843FF45082A801FF005155400FFD1420100055574AAA2AA800AA",
INIT_23 => X"AAA2D5421FF00042ABEFFF8400010082EAABFF55002ABEF087BE8ABA555168B5",
INIT_24 => X"E105D7BD7545A284020BA007FFFE10A284000AA0055401550055574005D2E800",
INIT_25 => X"0000000000000000000000000000000000000000000028B550051574005D7FFF",
INIT_26 => X"955455D556DA004971C7038140012482550E021C7EB8028A821C7BC516DFF800",
INIT_27 => X"17FF45E3DF471C70851400BA0071C5028FFD17FF6DAADB504001C71EDA82AAA0",
INIT_28 => X"FBE8B555D516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBF1D5492BED",
INIT_29 => X"C55554AAAAA480082FF84000BAEBF1FFF7DEB8000092552ABFFEF08517DF6DB6",
INIT_2A => X"087FEFA8241516DB55A2FFEAB6DEB843DF551C20801C71C5157428FFDB420101",
INIT_2B => X"5085550428412A85082BEDF401D71C0A2DBC7EB80000280824ADBD7490E28BEF",
INIT_2C => X"7D0051504005D71F8E004975D556DB68405092087FF8E00BE8A02082005F4714",
INIT_2D => X"A00557BD75EFF78000000000000000000000000000000000000000000000E2AB",
INIT_2E => X"200055557DE00A2801554555557FE100055554BA5504000105D2A80145AA842A",
INIT_2F => X"D7545AAD557410F7D57DF55AAFBD55450055420BA0055574BAF7D17DFFFAAFFC",
INIT_30 => X"ABDFFF08517FFFFF7FBEAB455D517FE00082EBDF45AA8428A10085568ABAA2FB",
INIT_31 => X"51554AAFFFFC00105D55554BAA28400000F784020BAAAD57FFEFA28402010552",
INIT_32 => X"8003FF55002AA8BEF007FFDE1000557DF45AAFBE8BEFA2803FF4555040015555",
INIT_33 => X"F7AE80000087BD55450855400BA002A95400F7FBC01555D2EBFF55A284000AA0",
INIT_34 => X"0000000000002EAABFF0051400105D5568A000051575FFF78415410087FEAA10",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000006000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"0202115002BB10080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"2FE962000017102918900948514522CE09200C0D590569398ADBF8CC1E50E480",
INIT_05 => X"5E6023002834854AE41C1E8782F508F2A15B71D412E0AFD9C2990DA56FF0B55A",
INIT_06 => X"82A803B9B9E55402000340003200220A86012D0000000480D02A7960540180A0",
INIT_07 => X"01380C40D890101DBD400901442800817C2901F400868554DE240000A80090CE",
INIT_08 => X"18A9050122004000005665510320C9C90510025A8A00000A0A048F550A440E00",
INIT_09 => X"2A8A562060410280081116C8204D016CB2CB2900080082795804112890000001",
INIT_0A => X"4052E400008176802200020025699200140001A15000017F0051D0F837324E00",
INIT_0B => X"5514554485D000000124002400000000000001004010A8812831605DA0000A05",
INIT_0C => X"708E2CB5320018CAC99BA0A3B9320018CAAAADA0C343F1AC1B01040A00202489",
INIT_0D => X"E7A3EE59320018CAC99BA0ACB9320018CAAAADA0CC421CA003B694B68018FAAA",
INIT_0E => X"24352AB2449A3FF2FA04E5E09B128834ADB1443A1891E4A928C29020E6A8524C",
INIT_0F => X"714C902375B801324301AB0067622E5E5404B2A5A40B1E6644AF0F021EA003AC",
INIT_10 => X"1216F50A8C241815FEB6A9158863F638FB60ED838E890B703C6260D8E3A21275",
INIT_11 => X"555E4C15F11133D171727A2550EE2F1BA0064F70DBDB1C74424E91E1C194C71D",
INIT_12 => X"ACCC59432A2B2D001F803471A9A960E57245FDF9D364DBD9435A6D45C9E81BED",
INIT_13 => X"0012CAC00006B0800000038814B72AB01508150013F162119014204373517700",
INIT_14 => X"002912300208092B940192D1000000000000A8A5AA80018120E0006600000000",
INIT_15 => X"1100011000110001100011000108000880008000520228080108039501200848",
INIT_16 => X"012000081500008A422150884081AC9000010003561180063DB4F61100011000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"28A28A3D2DE5F87963445469E79E7853D44C690DA64C1C69818768A360400000",
INIT_1B => X"F4FA3D3E8F4FA3D3E9A29A29A29A29A29A29A29A29A29A29A29A29A28A28A28A",
INIT_1C => X"000FA7D3E9F4FA7D1E8F47A3D1E8F47A3D1E8F4FA7D3E9F4FA7D3E9F4FA7D3E8",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"43FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE005500000000000000000000",
INIT_1F => X"80020005D2A95410FFFFC00000804154AA5D00001EFF78428AAA007BC2145F78",
INIT_20 => X"AD157400007BEAAAAAAAE955555D5568A105D2E974BAF7FBEAB45FFFFC00BAF7",
INIT_21 => X"007FC2000F78000010552E800AA002E821FFA2AAAAA00000417555FFD17DF45A",
INIT_22 => X"A08043FEBA5D55575FFF7AABFE00557BD74AAAAD17DF45F7D1421EF0055400AA",
INIT_23 => X"10FFD56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7AABDF55F7AE820A",
INIT_24 => X"FEF08517DF55A2FBEAB555D04154BAA2FBE8B55FFFFD55FF557FC2000FF80154",
INIT_25 => X"0000000000000000000000000000000000000000007FFDF45FF84000BA552ABD",
INIT_26 => X"28A821C7BC516DFF8438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE1049000",
INIT_27 => X"BE8B55FFF1C70BAF78A000005D2097438FFF1C7038140012482550E021C7EB80",
INIT_28 => X"0E1757DEBD17FF6DAADB504001C71EDA82AAA0955455D556DA00492490492F7F",
INIT_29 => X"3DF471C70851400BA0071C5028FF84020285D2085092002A801FFB6AAA8A1008",
INIT_2A => X"EBA4BAF6DE3AA8709208043FEBA555B555FFE3AABFE005D71D5492BED17FF45E",
INIT_2B => X"7557BC0028E38412428EBD16DA82410A3FFD7AAA4B8E824971F8E38E3DF45155",
INIT_2C => X"7DEB8000092552ABFFEF08517DF6DB6FBE8B555D04124BAB6FBE8B45E3FBD55D",
INIT_2D => X"55555003DE000000000000000000000000000000000000000000000000071FFF",
INIT_2E => X"00105D2A80145AA842AA00557BD75EFF78428B55AAD168B55F7FFFDFEFFFAA95",
INIT_2F => X"7FE10000000010F7FBEAB45FFD1554AAFFAE820105500154AAF7D5554BA55040",
INIT_30 => X"E801EFF7AEA8A10002E955FFA2D17DFFFAAFFC200055557DE00A280155455555",
INIT_31 => X"5557410F7D57DF55AAFBD55450055420BA0055574BAF784000BA5D0017410082",
INIT_32 => X"85568ABAA2FBD7545AA802ABEFA2AA9541000003DEBA557BD75EFA2AEBDE105D",
INIT_33 => X"FFFBEAB45AAFFD55555D7FC20AAA280000AAAAD17FE00082EBDF45AA8428A100",
INIT_34 => X"000000000000557FFEFA28402010552ABDFFF08517FFFFF7FBEAB455D04020AA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000002000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"5295B6957FCBE0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"6DE90201BF90102103AF158E805428249851BFB2C106592088DBF8400A5055C2",
INIT_05 => X"3824BD7F80148D9E07100A8201ED01C1A19B68F40A807ED9C18114956FF081DB",
INIT_06 => X"ED08CA6A8F033DD800000000050716BE9F57F8AC000807DFD999E0E5E1818B1B",
INIT_07 => X"00150886481240FE05A109228E2C0891D772A6F40045B8CF30E085DD2ED57D4E",
INIT_08 => X"72637FDF23800005981C0338190549C904182B6113870022000488C08B46268A",
INIT_09 => X"3E7437823DF78CDB6CA60E0E28EFFE2061872F80C1684A80C8604085F0074D3B",
INIT_0A => X"F5B4FFBD2FAD7FE653C36A1FF33E0E001E000B3A5DAADAFDDA5DA79350CFB801",
INIT_0B => X"CFE833C5C3D00018006C681700000000000000020012E9E10A31EB5FF9296A67",
INIT_0C => X"0D5ECE542A6FEEB2533EA160782A6FEEB2333EA16031F2BD47BDA2CA5D8164FC",
INIT_0D => X"282400F82A6FEEB2533EA160782A6FEEB2333EA160391BEFF2C32FB695F91911",
INIT_0E => X"573FAD5A86840354D1706FFFA3EF6E24B6D18C0D06638A207CFDE1F7DDAD76D5",
INIT_0F => X"FE4ACA4D77FAAB77CE3AF3EE78F58DB737E6E43E59AFE4A59B57679D19EFF2C7",
INIT_10 => X"ADB55572CA52606DFED6CA55334C04C04FF7D7A0ABD6DAAAB96529382B74E4E1",
INIT_11 => X"F9956EAA1A184045D5D7A870D2F5A5D7522D1281017F056E9C9C3FC95949C157",
INIT_12 => X"1F432EA58949D5B5C85F97871876F7D7E859FDEB974F486905001FDF5FA0D719",
INIT_13 => X"DEF20670021EE341036BF368128419FB5560158015177F916A039EF41FDB34A9",
INIT_14 => X"00633F1D0A7CC9AE7A08BFF0001D35682AC0CE8FCCC200A59BDD2FFE3F3EC7C7",
INIT_15 => X"FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A7800617112E46F05D02DD814102F8",
INIT_16 => X"05F08000179C16DECF67F08BC02F9086000D9E8A3F06ABD73DBCF4FBCF4FBCF4",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"34D34D48C4986868DC800181D75D7445F009EDCC4052E92E0204114F981800C0",
INIT_1B => X"1A8D468341A8D46834D35D74D34D35D74D35D74D34D35D74D35D74D34D34D34D",
INIT_1C => X"0008D46A351A8D46A351A8D46A351A8D46A351A0D068341A0D068341A0D06834",
INIT_1D => X"0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"43FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF5500000000000000000000",
INIT_1F => X"8028A00F7843FEBA55043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE00550",
INIT_20 => X"804154AA5D00001EFF78428AAA007BC2145F7D568B45000002010552EBDF45A2",
INIT_21 => X"5D2A95410FFAE800105D2A95410002A95410AAAEBFF55AAFFC00BAF7FFC00000",
INIT_22 => X"FFFD57DE00F7AE800AAAAAABDFEF5D2E974BAF7FBEAB45FFFFC00BAF78002000",
INIT_23 => X"AA5D517DF45AAD157400007BEAAAAAAAE955555D5568A105D7FFFFEFA2D568BF",
INIT_24 => X"1FFA2AAAAA00000417555FF8028B55082A974105D003FF55F7802AAAAAAD168A",
INIT_25 => X"0000000000000000000000000000000000000000000000010552E800AA002E82",
INIT_26 => X"955C71C043FE10490A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD749000",
INIT_27 => X"E050384124BFF7DB68A28A38F7803DE82490438FC7E3F1EAB55B6DF6DBFFF7AA",
INIT_28 => X"F5C70BAFFF1C7038140012482550E021C7EB8028A821C7BC516DFFDF68B551C0",
INIT_29 => X"FF1C70BAF78A000005D2097438FFAA85000492495428082E95400AAA0BDF7DB6",
INIT_2A => X"497FFAFFFB6D56FBFFEBDB78E38F7AA800BAB6AEBDFD75D2490492F7FBE8B55F",
INIT_2B => X"DEB8028AAAB6D16FA8249517FF6DAADB504001C71EDA82AAA0955455D556DA00",
INIT_2C => X"285D2085092002A801FFB6AAA8A10080E1757DEB8A2DB5514249243841003FF6",
INIT_2D => X"0BAF7FFFDF550000000000000000000000000000000000000000000000004020",
INIT_2E => X"8B55F7FFFDFEFFFAA9555555003DE00002ABFFEFF7FBFDFFFAAD168B55AA8000",
INIT_2F => X"D75EFF7FBEAB45552E954BA08003DFFFFFAAA8AAAF7843FE10000428B55AAD16",
INIT_30 => X"E95410AA843FFFFF7D5554BAF7D5554BA5504000105D2A80145AA842AA00557B",
INIT_31 => X"0000010F7FBEAB45FFD1554AAFFAE820105500154AAF7AE974000800154AA002",
INIT_32 => X"2801554555557FE10007FEABEFFFD57FFEFAAFFE8ABAFFAA820BAF7AEBFF5555",
INIT_33 => X"5500020AA08003DFFFA28028AAAF7D17DE0000517DFFFAAFFC200055557DE00A",
INIT_34 => X"00000000000004000BA5D0017410082E801EFF7AEA8A10002E955FFA2AABFF45",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000067FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"080BA868803F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"42016B0C401F58495C900A4859552A611D9A640F5903B2388004004C08A06008",
INIT_05 => X"16226B107811422A641C08038040007060E0032801E0202000991B708280B501",
INIT_06 => X"120886B3B8E0FC86142B4142B0000000011114D3058240240907F82000000000",
INIT_07 => X"006880802102401015610A02C4005000EA019D002482043FCF1C8090C02800C0",
INIT_08 => X"11018020D40A5004003260F9810541494D403D9B98810A0002C601000054B94A",
INIT_09 => X"022E0C6070000504102805C820C8016C30C250080C0182183804012A0A102200",
INIT_0A => X"084001E000108010230495A800FD865421432121804021C20452880C2D100000",
INIT_0B => X"3F140FC2060014250B9080008306C18360C1B0609C05013065CC042004040808",
INIT_0C => X"DF7C728582081483ACC15F9C3982081483CCC15F9CBA45505640000A40201900",
INIT_0D => X"DFEBFBF982081483ACC15F9F3982081483CCC15F9FB1962FCB69E08AAAEAEBCD",
INIT_0E => X"CAA02FE3F8E7F5E3AC3620805298B15A3FEBF1CFFF7670ACC3811A28AB57523C",
INIT_0F => X"01BD67DC4041D4CF03138DD865103EFEEAC9002BF05800D875E63CC9962FCB52",
INIT_10 => X"0016EA8DB7BFE25208E8F46A228BF8A757F1B72A8A800B7546DB9F1CA320037F",
INIT_11 => X"81A8A29509EAAE7FD3B749471C48F8A45981CCFAFDBF9464006FD037AEFAE515",
INIT_12 => X"EFF5778802A3AF8E8FB0440CE78773B709641256EC844B8AF92FD7CEDC24A9E1",
INIT_13 => X"0003C1C284601C2864000080113307E4800297D086E00036D2440E0880AAD62B",
INIT_14 => X"C44C92A88DCC2211E44174112840880000060D7030C30B885200D27400400808",
INIT_15 => X"0030800308003080030800308001840018400400602A01880980037109700C04",
INIT_16 => X"6808348340000020301805002D008CD943626111C0D95C20C2030A0030800308",
INIT_17 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B0",
INIT_18 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_19 => X"00000000000000000041B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_1A => X"1451451223059150A2EFB05C104104B3CEB80EE173C2300FCA8B7DF160000000",
INIT_1B => X"4AA552A954A25128955545145145155555545145145155555545145145145145",
INIT_1C => X"00025128944A25128944A25128944A25128944A25128944A25128944A2512894",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"43FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA0000000000000000000000",
INIT_1F => X"8400145AA801741000043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF550",
INIT_20 => X"7FBE8B45AAD568BFFFFAA975FF00003FE0055043FFFFFFFFFDFEFA2D56AB45AA",
INIT_21 => X"F7843FEBA55557FFEFA2D168B55AAFBFFFFFFF80021EF0855421EF00043FFFFF",
INIT_22 => X"A5D2A82155F7AEBFEBAFFD56AA00A2D568B45000002010552EBDF45A28028A00",
INIT_23 => X"BAA2FFC00000804154AA5D00001EFF78428AAA007BC2145F7D5400000004020A",
INIT_24 => X"410AAAEBFF55AAFFC00BAF7AE80010082E954BA0004174AAAA8428B45082ABFE",
INIT_25 => X"0000000000000000000000000000000000000000002E800105D2A95410002A95",
INIT_26 => X"00038F7DB6FBD7490E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA55041549214000",
INIT_27 => X"1F8FD7AAD16FB6DBE8E00155BE8015410140A3FFFFFFFFFDFEFE3F5FAF45AA80",
INIT_28 => X"5B471C7140438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE1049043FFEFE3F",
INIT_29 => X"124BFF7DB68A28A38F7803DE82495B78FC7AAD56FB6DBEF1FAFD7E384001EF14",
INIT_2A => X"FFD1420381C0A02082492A85155E3A4BDE92FFD56FA28B6DF68B551C0E050384",
INIT_2B => X"ABE8E28B7D1420BDEAAA2F1C7038140012482550E021C7EB8028A821C7BC516D",
INIT_2C => X"00492495428082E95400AAA0BDF7DB6F5C70BAFFAE870280024904BA1400174A",
INIT_2D => X"4BA550415410550000000000000000000000000000000000000000000002A850",
INIT_2E => X"DFFFAAD168B55AA80000BAF7FFFDF55002ABFFFFFFFFFFFEFF7FBFDFFFF7AA97",
INIT_2F => X"3DE0000043DFEFA2D56AB45AAD57DFEFF7AA82155F78015400552ABFFEFF7FBF",
INIT_30 => X"568B55A280021EF557FD7555550428B55AAD168B55F7FFFDFEFFFAA955555500",
INIT_31 => X"FBEAB45552E954BA08003DFFFFFAAA8AAAF7843FE10007FEAB55A2D17FFEFFFD",
INIT_32 => X"A842AA00557BD75EFF7D1400AA5D2A82000002A95545A2843FE00F7D17FEAAF7",
INIT_33 => X"0004020AA5D04154BAF7AEA8BEF55003DEAAA2D5554BA5504000105D2A80145A",
INIT_34 => X"0000000000002E974000800154AA002E95410AA843FFFFF7D5554BAF7AE974BA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000002000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000010228001000000000000000000024001620280000000000354200004008",
INIT_04 => X"00016200001310090090004840004152C7208802590000388000004C08006000",
INIT_05 => X"1621008008100002641C0803804000702000000000E02000009900000000B100",
INIT_06 => X"00A0010210200C00000000000000000000000080000000000000D82000000000",
INIT_07 => X"010084C00D267001B880080700285020020AC988200228024004804050089011",
INIT_08 => X"0E0E00000000000000106009872048400C4000010D000008000204150A00815A",
INIT_09 => X"022A040000000000000004C80000002C30C20000000002180800580000000000",
INIT_0A => X"0007600000000000000000080025860000000080A00020602040800000000000",
INIT_0B => X"031400C002000000000000000000000000000000000000000000000000000084",
INIT_0C => X"28DC0D385598035D0008A003B05598035D0008A0034078104B41A41000000000",
INIT_0D => X"041124505598035D0008A000B05598035D0008A0004263C0343EDD4140040422",
INIT_0E => X"B740500401180DE053A98F6ECC739D8140040231068187C39F5A4F985C008902",
INIT_0F => X"000010227848D4303807FC8CC5508AEAED1BFBD406451B02000E033263C0343C",
INIT_10 => X"D6480000000018A700FCF980CC300318A2420851546B2400000040D8549B5800",
INIT_11 => X"81C21140E40511802208D6B30C48F8A8A452210402120A936B0000000004C2A8",
INIT_12 => X"F9E9410006362A2B6424287B08286208D6B1427ED430B41402D0250823597001",
INIT_13 => X"0002C040000000000000000010030060009C000018440021011821B35254E99A",
INIT_14 => X"000040002000044000000000000000000002F0001F00002024B2000200000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"00000000000000000000000000008C8000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C30C30D0A208C4DC822EC1534D34C01FA3F0C7010C6600A0200441920000000",
INIT_1B => X"26130984C26130984C30C30C30D34C30C30C30C30D34C30C30C30C30C30C30C3",
INIT_1C => X"000130984C26130984C26130984C26130984C26130984C26130984C261309A4D",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D00000000000000000000",
INIT_1F => X"AA974BA5D517FFFF08043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA007",
INIT_20 => X"FFFFFFFFF7FBFDF55A28402000F7D56ABFF557BFFFFFFFFFFFFFFFFFBFDFEFFF",
INIT_21 => X"AA8017410007BFFFFFFFFFFFFEFF7D16AB45AA8002000F7D5575455D043FFFFF",
INIT_22 => X"5AAD568B55F7AE955FFAA840201008043FFFFFFFFFDFEFA2D56AB45AA8400145",
INIT_23 => X"FF5D043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE00557BFFFFFFFFBFDF4",
INIT_24 => X"FFFFF80021EF0855421EF002ABFFEFF7D168B55AAD17FFEFF7AE975FF00557FF",
INIT_25 => X"000000000000000000000000000000000000000000557FFEFA2D168B55AAFBFF",
INIT_26 => X"954AA5504154921471FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA55000008255000",
INIT_27 => X"FFFFEFF7FBFAFD7E3A4954BA555B7AFC7080E3FFFFFFFFFFFFFFFFBFDFEFFFAE",
INIT_28 => X"DF52545550A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD74975FFFFFFFF",
INIT_29 => X"AD16FB6DBE8E00155BE8015410147FFFFFFF7FBF8FC7EBD568B55A28000000FF",
INIT_2A => X"497BFDFC7E3F1FAF55A2DB6FB7DF7AE955C7BE800000008043FFEFE3F1F8FD7A",
INIT_2B => X"7EBA0955FF145B7AFC7410438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10",
INIT_2C => X"C7AAD56FB6DBEF1FAFD7E384001EF145B471C71424B8FC7E3D56AB6DB6DF7AFC",
INIT_2D => X"4AA550002000550000000000000000000000000000000000000000000005B78F",
INIT_2E => X"FFEFF7FBFDFFFF7AA974BA55041541055517FFFFFFFFFFFFFFFFFFFFEFF7AA97",
INIT_2F => X"FDF5500517FFFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB45002ABFFFFFFFFF",
INIT_30 => X"56AB55A28002000F7FFC2155552ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FF",
INIT_31 => X"043DFEFA2D56AB45AAD57DFEFF7AA82155F78015400557BFDFEFF7FBEAB55A2D",
INIT_32 => X"FAA9555555003DE00007FFDF45AAD568B45AAFBFFFFFFFAA95545F7840201000",
INIT_33 => X"AAD16ABFFFFFBEAB45A280155EF557FE8B55000428B55AAD168B55F7FFFDFEFF",
INIT_34 => X"0000000000007FEAB55A2D17FFEFFFD568B55A280021EF557FD755555042AB55",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000004000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"0001E6000053300B00D0005800000000000000407B0004BB830004DC3D01E000",
INIT_05 => X"FEE0000008720043EC3C3D0F87FA19F7E0201C409BE1F10623BB000A100CF300",
INIT_06 => X"00200006102FFC8E0007C00078008000171175A200096404D97FFBE4744200AA",
INIT_07 => X"000000482491301000010001DC00000000000000004203FE4005800000008030",
INIT_08 => X"40800020E2008000027FEFF946058180010429000001080AAA010F8000000000",
INIT_09 => X"03EAFE400000120000913FD80000003DF7DE0080010047FBF8000000000800C5",
INIT_0A => X"0800000080000010000400080FFDBE0000004000000100000100506002204610",
INIT_0B => X"FF14FFC00600000000801020000000000000010240001721214E000004000000",
INIT_0C => X"A70C0008020000200000000F30020000200000000F3008001E00000000001803",
INIT_0D => X"004A58F0020000200000000F30020000200000000F3040200000020000000026",
INIT_0E => X"000000000019B140000800800000020000000030B86000400080000200000000",
INIT_0F => X"000014AC08000000508001030A0A4001000000000002183E61E6000040200001",
INIT_10 => X"0000000000A56000090100000000001F86C00010080000000000525801000000",
INIT_11 => X"0600000000001716800000803102020000000002BC360020000000000292C010",
INIT_12 => X"06049CDF70C08040100000706707600000801000000000000057450000100106",
INIT_13 => X"000ADFC011001C81080001101F977FE008000000000000400400400020000805",
INIT_14 => X"0000000000000000000000020020029000000000000000020000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000002000200000000",
INIT_16 => X"0080800801810100000000000093ED8000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000401",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"18618640C49821201C0001A1E79E79A4B0038200010089054C1A0104D2040020",
INIT_1B => X"0C86432190C86432196596596596596596596596596596596596596586186186",
INIT_1C => X"00086432190C86432190C86432190C86432190C86432190C86432190C8643219",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA5504020100800000000000000000000",
INIT_1F => X"AA974AA550002000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7",
INIT_20 => X"FFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFFFFFFFFF7",
INIT_21 => X"5D517FFFF087FFFFFFFFFFFFFFFFFFFFDFEFFFAE974AA5D003FE005D043FFFFF",
INIT_22 => X"FF7FBFDFFFAA84000105D556AB55557BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA",
INIT_23 => X"EF08043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55003FFFFFFFFFFFF",
INIT_24 => X"B45AA8002000F7D5575455D2EBFFFFFFFFFFFEFF7FBEAB55A28000010F7D16AB",
INIT_25 => X"0000000000000000000000000000000000000000007BFFFFFFFFFFFFEFF7D16A",
INIT_26 => X"954BA550000082557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA55040002800000",
INIT_27 => X"FFFFFFFFFFFDFEFF7AE974BA5500050380071FFFFFFFFFFFFFFFFFFFFFFFF7AA",
INIT_28 => X"0038E285D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA55041549214043FFFFFFF",
INIT_29 => X"7FBFAFD7E3A4954BA555B7AFC70871FFFFFFFFFFFFFFF7FBFDFFFFFAA974BA55",
INIT_2A => X"490E3FFFFFFFFFDFEFF7F1FAFC7A28002028555F6FB7D5D75FFFFFFFFFFFFEFF",
INIT_2B => X"5A28402010FFDB6ABEF140A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7",
INIT_2C => X"FFF7FBF8FC7EBD568B55A28000000FFDF525455524BFFFFFFFBFDFC7E3F5E8B4",
INIT_2D => X"4AA5504000BA080000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFEFF7AA974AA550002000557FFFFFFFFFFFFFFFFFFFFFFFFFFAE95",
INIT_2F => X"1541055043FFFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08517FFFFFFFFF",
INIT_30 => X"FFFFEFF7AE974AA550028AAA5D2ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA5504",
INIT_31 => X"517FFFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB4500557FFFFFFFFFDFEFF7F",
INIT_32 => X"A80000BAF7FFFDF55002EBFFFFF7FBFDFEFFFD568B55A284020BA557FFFFFF5D",
INIT_33 => X"F7FBFFF55A2D16AB45AA8402000F7FBEABEF5D2ABFFEFF7FBFDFFFAAD168B55A",
INIT_34 => X"0000000000007BFDFEFF7FBEAB55A2D56AB55A28002000F7FFC215555043DFEF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"1094EC681244819000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"0001E6000053300F01D4587800446194F49020107F0012BBC00202DC3823EA82",
INIT_05 => X"FFF201B228704123FC3C381F87C03DFFF012412A9FE1E01013BF09404050F300",
INIT_06 => X"100B3096F43FFF002004020044041084CB01AD0000037617027FFFE050000080",
INIT_07 => X"A12034043C802A821D41412001A0040950AB60014114C3FE4187A009A663A680",
INIT_08 => X"7F40002C01004000047EFFF811A46968004060629A0002208A00000068113205",
INIT_09 => X"E3EBFE0A812D8D5B742D3FF84056383FF7DE0880042107BFF9C45B85101C49A3",
INIT_0A => X"02804A08221890004806C0310FFDFE00040009814C089202225412115414601D",
INIT_0B => X"FF56FFC0281280080180B2948004400220011100841200D001000624000100C0",
INIT_0C => X"50025360694101816002D41A4068C101815004D8158809C86065941840B1014F",
INIT_0D => X"82418A0068C101816002D41A40694101815004D815810D42E04A08A80098C024",
INIT_0E => X"1A300012682960828F05C96A001B029010134160C8125B0B271802242880A044",
INIT_0F => X"49F115100920C54E8EA256ECF078BA081C10080E05C0B06AA8B12CFD0D42E044",
INIT_10 => X"5144104F30A8801406D00290006280320100010362A8A20826A88660D86B2020",
INIT_11 => X"8010602011819E290048A2118EC8140C08064802C0081B0D64040936443306C5",
INIT_12 => X"C322A4C40A0300600C0A80509F418008804581BA0038005A706680012280506A",
INIT_13 => X"18DBFFC000120080002341881F3FFFF80DCC158092C044600466208CC5091011",
INIT_14 => X"806520398C6021569249C4B3007127080806FF917FC30010107688862A28C545",
INIT_15 => X"9228D9228D9228D9228D9228D99146C9146C84006309044081A001B188300E20",
INIT_16 => X"0448008004000000E07008010003EF80022A51904595123203040D9228D9228D",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_19 => X"0000000000000000004010040100401004010040100401004010040100401004",
INIT_1A => X"7DF7DF7FEFFDFDFFFBE7F3FCF3CF3FFF6EFF7FFDF7FF3EFC1FBFFDF7E0000000",
INIT_1B => X"FEFF7FBFDFEFF7FBFDF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF",
INIT_1C => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFD",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D00020000800000000000000000000",
INIT_1F => X"AE954AA5D00020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"55000200000003FFFFFFFFFFFFFFFFFFFFFFF7AA974BA5D0402000557BFFFFFF",
INIT_22 => X"FFFFFFFFEFF7AE974BA5D00174BA00003FFFFFFFFFFFFFFFFFFFFFFF7AA974AA",
INIT_23 => X"BA5D043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFF",
INIT_24 => X"FEFFFAE974AA5D003FE005D2EBFFFFFFFFFFFFFFFFFFDFEFF7AE954AA5500174",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFD",
INIT_26 => X"974AA550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000001000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"04050005571FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082557BFFFFFFFF",
INIT_29 => X"FFFFDFEFF7AE974BA55000503800003FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D",
INIT_2A => X"140E3FFFFFFFFFFFFFFFFFFDFEFF7AE954BA5D00154AA00043FFFFFFFFFFFFFF",
INIT_2B => X"FFFAA974BA5D00104925D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492",
INIT_2C => X"FFFFFFFFFFFF7FBFDFFFFFAA974BA550038E285D2ABFFFFFFFFFFFFFFFFBFDFE",
INIT_2D => X"4BA5D00000100000000000000000000000000000000000000000000000071FFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02000557BFFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7FFFFFFFFFFF",
INIT_30 => X"BFDFEFF7AE954AA5D041740055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5500",
INIT_31 => X"043FFFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08043FFFFFFFFFFFFFFFF",
INIT_32 => X"7AA974BA550415410552ABFFFFFFFFFFFFFF7FBFDFFFFFAA974AA5D00174BA08",
INIT_33 => X"FFFFFDFEFF7FBFFFFFF7AE954BA5D0000010552ABFFFFFFFFFFFEFF7FBFDFFFF",
INIT_34 => X"000000000000557FFFFFFFFFDFEFF7FFFFFEFF7AE974AA550028AAA5D2EBFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"8632CA211E4491D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"24B000808800040439245B221373581F97B0A8D1040F92000F42000047A00E58",
INIT_05 => X"011B2BBA308F023810004700083E220811E9BF2844021B1004045E4249500449",
INIT_06 => X"EF018980A51003AA0200C020088E16A85235722940A817251100040D6D0702A2",
INIT_07 => X"24E8145C9ECAB0D247B013B405EAD525FAE48FC2060B880081A26DCD4047EFF9",
INIT_08 => X"0050482D0141C0055280100751096B6A40D6F86723E510AA2004803D3275EB20",
INIT_09 => X"20110204804818CD280100207246A8020000AC0283002004051507A5411C0DA0",
INIT_0A => X"4E506A2C6898B2950AA6D635B00041C23020131A80CFDFF3FE509A907C556828",
INIT_0B => X"002200050F60E220A06880D2A14050A028501428054278142151262CA5034385",
INIT_0C => X"F06273612B3482C0C0078E1F412B1582C090078E1F840A2B0114020104022460",
INIT_0D => X"C2C0DB012B1582C0C0078E1F412B3482C090078E1F891C239F8908003099C1AC",
INIT_0E => X"0828041BA859F213AFC14AA380430060181BA1B0FD16770236A4091621C08055",
INIT_0F => X"095337B08AA600CA88B143AB11880C280600101F09C030AB28B03C111C239F87",
INIT_10 => X"3096004B61BD8068B92400D0004E30368910E8822A984B0025B0DE6089462660",
INIT_11 => X"F07830001AC2173B00E162563454C40804055412D4481128C4CC012A66F30455",
INIT_12 => X"BF006850840180A00E1C81900C4190E160589C48082C006A9057CA4385809520",
INIT_13 => X"39C020004416B105036B4180C000800C8C00460848952220592745AC11A544B1",
INIT_14 => X"103D2A512C6A8C4F0008AA800470370000A0004D0000002126F30C902A29C545",
INIT_15 => X"C2A81C2A81C2A81C2A81C2A81C9540E1540E001400006100003202D040050220",
INIT_16 => X"45E22022365034A8EA754008004C0214202C50013456520CA09281C2A81C2A81",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"0040100401004010040100401004010040100401004411044110441104411044",
INIT_19 => X"0000000003FFFFFFFF9004010040100401004010040100401004010040100401",
INIT_1A => X"3CF3CF7FE7FDFD7DF7EFFDDDF7DF7DF7DEFE8FF1F7DEBD6FCD9F7DF7D0512289",
INIT_1B => X"FE7F3F9FCFE7F3F9FCF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"0007F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04000000000000000000000000000",
INIT_1F => X"AE974BA550000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D00020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00000AA007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAA954BA5504000AA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA",
INIT_23 => X"BA5D7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFF",
INIT_24 => X"FFFF7AA974BA5D040200055517FFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500000",
INIT_25 => X"000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040200008000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"00020BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D",
INIT_2A => X"5571FFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5504020AA5D7BFFFFFFFFFFFFFFF",
INIT_2B => X"FF7AA974AA5D00070925D71FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082",
INIT_2C => X"FFFFFFFFFFFFFFFFFFEFF7AA974AA5D040500055517FFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D040200008000000000000000000000000000000000000000000000003FF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAA954AA5D00020AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504",
INIT_31 => X"7BFFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7BFFFFFFFFFFFFFFFFF",
INIT_32 => X"7AA974AA55000200055517FFFFFFFFFFFFFFFFFFFFEFF7AA974BA5504020BA55",
INIT_33 => X"FFFFFFFFFFFFFFDFEFF7AE974AA5D00154105D517FFFFFFFFFFFFFFFFFFFFEFF",
INIT_34 => X"000000000000043FFFFFFFFFFFFFFFFBFDFEFF7AE954AA5D041740055557FFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"5886C0201A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"0005EE040057700F40D08078500000D9218020407F0000BB8018A2FC380BEAC2",
INIT_05 => X"FFE0419028700023FCBC385F87C0BFFFE0124002FFE1E0C517FF09111212F300",
INIT_06 => X"DF0AF116D03FFC96102081020000020489019C4304802412027FFFE000000000",
INIT_07 => X"B710000001160A003475C8100123400E20E1F40F439647FF4807E189A477EF81",
INIT_08 => X"7F0F94801008000007FEFFFB110140695812CC4188D58A0AAA10803448D0844F",
INIT_09 => X"C3EBFD4201258112D4487FF8001010FFF7DE4000000003BFF8C2581808002001",
INIT_0A => X"0801000C024000004A9400000FFDFF50010103134CAFDF03BA18000F39900037",
INIT_0B => X"FF57FFC02812F00429DC92C40002000100008000105400C00400100000A01800",
INIT_0C => X"424202A1CAF13F214001521001CBF03F21100152100801C17E61841950B1C10F",
INIT_0D => X"420B8001CBF03F214001521001CAF13F2110015210088528E00E02C8200A430A",
INIT_0E => X"12480202C86040902AC60BACDF0E02D02001C1C044006D0C94FB94320880603C",
INIT_0F => X"09B00300010AF5052419D196441902801430182800A018D9CA8000648528E00D",
INIT_10 => X"C140004D101808458A5602E000892029110445C19960A00026880C0067390000",
INIT_11 => X"4040301009408021144CB042F880100C0601844068880CE72000013600600332",
INIT_12 => X"EE38A1F80E02120018390320F050144CB241D0B9023402085020825132C8CB5B",
INIT_13 => X"001BFFC200400020224000405F7FFFE0008E17C0D240406519400500840A9524",
INIT_14 => X"907120AC810033149249C433200180082A06FF907FC308181204800600000000",
INIT_15 => X"1010C1010C1010C1010C1010C10086080860840063090442A18001B188300C48",
INIT_16 => X"2000100100000000000004002403EFC10302219A41C1443243050C1010C1010C",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_19 => X"0000000000000000000080200802008020080200802008020080200802008020",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"550000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974AA550400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"00087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE954AA5D00000AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA5504020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA55",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400010087FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE954AA5D0402038007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE954AA5D00020BA087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"00010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D00",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA55040001000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAA954AA5D04000AA087FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D00020AA007BFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"0000745C200801000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"0001E6000053300F00D0007810042140C00000407F0000BB800000DC3801EA00",
INIT_05 => X"FFE0000008700003FC3C380F87C019FFE01240009BE1E00003BF00000000F300",
INIT_06 => X"DC8C3006103FFC0000000000000000048900880100800012027FFFE000000000",
INIT_07 => X"0061200009B24B043980021000810284204A8001401643FE4007E5501AA00000",
INIT_08 => X"7F00000000000000007EFFFB11A56940581280031D61420000B080102040BC5B",
INIT_09 => X"C3EBFC020125811254083FF80000003FF7DE0000000003BFF800580000000001",
INIT_0A => X"0580000000000000000000000FFDFF4000000AA0354000019C40000128000011",
INIT_0B => X"FF56FFC000104000000010440000000000000000001000C00000000000000240",
INIT_0C => X"48C0804012500021B00880108012500021E00880104809C1666594584031010F",
INIT_0D => X"0501840012500021B00880108012500021E0088010492064206100E810842000",
INIT_0E => X"0270040410004C840041A0D8005410903804100144800803419043064900C002",
INIT_0F => X"400041020902F60002260D65B361BAA1041018140F02C0000809408D20642053",
INIT_10 => X"D0021800020818B06D9802F00030C02060110002C9E8010C00010480B35A0300",
INIT_11 => X"90203020042108603100061516EE800C060228204300166B4060080008240593",
INIT_12 => X"14AE4C7C02000040206602C10B48110006143B62023C00142800B04400095DFF",
INIT_13 => X"001BFFC000000000000000001F17FFE000DC1180C78044000440292083010402",
INIT_14 => X"814080008000010012414433000100080806FD107FC300000000000600000000",
INIT_15 => X"1000C1000C1000C1000C1000C100060800608400630104408180012188300C00",
INIT_16 => X"0000000000000000000000000003EF80020201904181003003000C1000C1000C",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"3DF3DF64C7986120B42BB99575D75FFD2AF6E7CC1132CD73DF3A441990000000",
INIT_1B => X"1E0F0783C1E0F0783DF7DF7DF7CF3CF3CF3CF3CF3DF7DF7DF7DF7DF7DF3DF3DF",
INIT_1C => X"0000F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100800000000000000000000",
INIT_1F => X"AE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"00007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D00020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010080000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000001008",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA550000010087FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002010087FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00004000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"4909E6093253306F82D0007C80000000080E01007F8020BBC00040DC3801EA00",
INIT_05 => X"FFE0000008704503FE3C380F87C019FFF01241009BE1E00203BF80800000F392",
INIT_06 => X"CC083006103FFF9E2086C2086E006604C9019D03108B7412027FFFE070400880",
INIT_07 => X"0000004024057000000100000000000000000001401643FE4007C00000000000",
INIT_08 => X"7F00000801404000007EFFFF40010000401408000045000000A0801000408000",
INIT_09 => X"C3EBFF4A7DF795965C6D3FFC0020003FF7DF01880C618FBFFDD75E0010004043",
INIT_0A => X"0000000000000000009400000FFDFFC006020000000000019804000028000191",
INIT_0B => X"FF56FFC02812E0182000F2C48304418220C11160845004D04820000000000000",
INIT_0C => X"0800800002400001000800000002400001000800000801C0786184185031810F",
INIT_0D => X"0400000002400001000800000002400001000800000000202000000800000000",
INIT_0E => X"0200000000000404000000880000001000000001000000000090000008000000",
INIT_0F => X"000040000100C600800001040000040009100000000200200000400000202000",
INIT_10 => X"4000000002000000081001000000000040010000082000000001000001080000",
INIT_11 => X"0000400080000040010000001080001008000000010000210000000008000010",
INIT_12 => X"0420000000030280000000010000010000001020000000000000100400000108",
INIT_13 => X"001BFFE0120012C1400080291F17FFF0018C11808200400000400000C2000000",
INIT_14 => X"80400000800001001243443B000100880806FD107FC301800000000600000000",
INIT_15 => X"1000C1000C1000C1000C1000C10006080060840077330C4889CC292588300C00",
INIT_16 => X"44C82082068C0200000008014023EF80020201904189003003000C1000C1000C",
INIT_17 => X"4110441104411044110441104411044110441104411044110441104411044510",
INIT_18 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_19 => X"2FFFFFFFFFFFFFFFFFC110441104411044110441104411044110441104411044",
INIT_1A => X"0924821409005312E8A25E15A69A6BFB0A196A8C5A2932F7C13C15DA08080000",
INIT_1B => X"C46231188C462311892492492492492492492492482082082082082082092482",
INIT_1C => X"00162B158AC562B158AC562B158AC562B158AC562B158AC562B158AC562B1188",
INIT_1D => X"0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"00087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04000",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040200000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"94A7B2B1450000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"6FEBEF5FEC737AFBC6F85FDEB220109E1FEFFFE3FBA7FDFB9BD301DC3FF5F0D2",
INIT_05 => X"FEEDBFDC387F987FEF7C3FAF87FF59F7F5FB7FF59BE1FF980BBBB7FE6D21F3DB",
INIT_06 => X"DFA08957902FFDEE9D7DC9D7DF2B263893479DDFAFDFE15213FFFBE1F1D3A333",
INIT_07 => X"00018010992310605CE10301DE0C1831CB7DF60A244B9BFEE00589DDBCEFEDC1",
INIT_08 => X"FFEFAA001D8EA111DA7FEFF90F21C8C84D9C0D858FC7020828C18FD18346BBF0",
INIT_09 => X"0BFAFFF37DF7B9DF7DCB3FDE89ECC07DF7DF5F985C6BCFFBFA28F99E7EB07F47",
INIT_0A => X"0607307DCFE1D4077B4D0026FFFFBE7D67D7F3BB79CFFB83BF14EC1E7D598058",
INIT_0B => X"FFFCFFC7D7D51D6F5FDCB935D7AFEBD7F5EBFBF7FEBD66DBFCA3F87501AE7B08",
INIT_0C => X"40520201F45EC0010007E01001F45EC0010007E010084BCD7FF1B61B5C33813F",
INIT_0D => X"0001A001F45EC0010007E01001F45EC0010007E01001BD8020500008001F0100",
INIT_0E => X"0200001EC00040B02007EC09A0E00010001DC0004600400F781429C008000077",
INIT_0F => X"81C203404B3BFD0402346235408402C08010003C064000E408010081BD802060",
INIT_10 => X"68B1000E401A08FE0012040000FC002001360403E434588007200D00F88C84C0",
INIT_11 => X"281D00001F01002156040675809145400007B00040091F1190982038406807C8",
INIT_12 => X"903A80008320C0403C34000088601604067D00212000007C400082D81009FC08",
INIT_13 => X"D6BFDFF7BFFED3FBFF6A84383F177FF005FFBFF5FA1040076065F730FC08043A",
INIT_14 => X"CDEBCFF589807B7096CD4CF73AC1FC98884FFF19FFC71FEFED7B251E35768E8E",
INIT_15 => X"78C0D78C0D78C0D78C0D78C0D7A606BC606B8C56F7730ECCDBDF152199F51EDD",
INIT_16 => X"FEFDFDDFE7DD87FEFF7FF796FFFFFDFFD7E681B867D3683A03A40F78C0D78C0D",
INIT_17 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFB",
INIT_18 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_19 => X"6FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_1A => X"4C30C375E2BD54D5D6C565F871C71D44FCF491E166CC853E8695F86EDB5C8864",
INIT_1B => X"26130984C26130984C30C30C30C30C30C30C30C30C30C30C30C30C30C30D34D3",
INIT_1C => X"000130984C26130984C26130984C26130984C26130984C26130984C26130984C",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"1085B0B041000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"6FAB975B6470BAF386C87A9CB00000001FEF9F23E3A7BDE79B5101D23FB5C0C2",
INIT_05 => X"F8EDBFD4347F18778E723F2E47FE59C7F5FB7F759B91FB880BA3B6FE2921CBDB",
INIT_06 => X"DFC00147000FFC128D5CE8D5CC210638A046889CAB57E84217FFE3E181932377",
INIT_07 => X"000141000000042000000288020C18300320620A80231BFE200181092CE7ED80",
INIT_08 => X"FEEF22000C562551D87E8FF90041101042110180004102800008801183468180",
INIT_09 => X"0BE0FC137FF7A0FF75813F1C85244071EFBF17D85C738BE3FA08F9DE36B05B07",
INIT_0A => X"040510768EA0C406630D00226FFE3E2D62D6E21259CFDB039E806C0245188040",
INIT_0B => X"FF48FFCC57550D63564D1D2556ADAB56D5AB6AD7EAB962CBD8A3A83101F47E08",
INIT_0C => X"00130201E44A40010007600005E44A4001000760000843C561E5C55C42B9011F",
INIT_0D => X"00002005E44A40010007600005E44A40010007600004BD8020100008001F0100",
INIT_0E => X"0200001EC00000382006EC0820A00010001DC0000208400D781020C008000077",
INIT_0F => X"81C20040431BC50402146235400400408010003C064000C400018080BD802020",
INIT_10 => X"4821000E400204FE0010040000FC0000003E0403A424108007200102E8888080",
INIT_11 => X"080500001F0100005E040475808101400007B00000015D111010203840081748",
INIT_12 => X"903A8000012040403C34000080201E04047D00202000007C400000F81001FC08",
INIT_13 => X"109E1FE5ADA4C25ADE72041A3F147FF0018DBBB5FA10400360649310FC08003A",
INIT_14 => X"EFABC7054880693016DD4C755AC16C1A884FFE18FFD757E7ED7A211E81C09818",
INIT_15 => X"3440C3440C3440C3440C3440C3C2061A2061AD46FF730E5CCBCD55219AB55F0D",
INIT_16 => X"DE75ED5EC71385FC2512E3565BBBF1BAD6F281BC63F1683803C00E3440C3440C",
INIT_17 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6B",
INIT_18 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_19 => X"7FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_1A => X"0000003C010072F24388521000000140A8100481CA8604368714104A47168874",
INIT_1B => X"8040201008040201000000000000000000000000000000000000000010400000",
INIT_1C => X"00140A05028140A05028140A05028140A05028140A05028140A05028140A0100",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"8C2100804900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"02000100440408002408008002221000204116A280000F000001400000100010",
INIT_05 => X"0004D44400004D4400000000000000000000005C0000000A0000002C20600000",
INIT_06 => X"2000004100000120040A0040A00B009000620294010000400080000888800911",
INIT_07 => X"2488045002489020420110800244891211440804000810002000081040000000",
INIT_08 => X"00B062080542C004CA00000050080202008401842004108AAAA00008912240A1",
INIT_09 => X"2800010000000C0000E400002040500000009202C10020400044000222000204",
INIT_0A => X"02043058C460540329810002D002000400407020800000004000640800088008",
INIT_0B => X"0008000140000401028008330000800040002002480102010082981500062108",
INIT_0C => X"00500000040A40000000A00000040A40000000A0000040060084104110828030",
INIT_0D => X"00012000040A40000000A00000040A40000000A0000000800010000000000000",
INIT_0E => X"00000000000000A00000040020A000000000000006000000080020C000000000",
INIT_0F => X"8000024040152000000020000004004080000000000000240000000000800020",
INIT_10 => X"0821000000120002000004000000000001220000040410800000090000808080",
INIT_11 => X"0805000000000001420000200001014000000000000900101010200000480008",
INIT_12 => X"0000000001204000000000000820020000200000200000000000028800002000",
INIT_13 => X"29400000933050080C0001900020000000408010000000022000D61028000008",
INIT_14 => X"440245400082D022040000400800081022C0000080000206CB0821082B694D4D",
INIT_15 => X"605016050160501605016050160280B0280B0012000843066021001400040024",
INIT_16 => X"0810840861CD33548542A10209D4100E4040A00002002C004001036050160501",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008021",
INIT_18 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_19 => X"0000000000000000000020080200802008020080200802008020080200802008",
INIT_1A => X"41041001A835050788440B58C30C31DF6C110A00246972C0C39989A40A0C22E1",
INIT_1B => X"C06030180C060301810410410410410410410410410410410410410410410410",
INIT_1C => X"00160B0582C160B0582C160B0582C160B0582C160B0582C160B0582C160B0180",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0803B2814D0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"26E1E905CC574828C4F85FC600000016004F77E2F887CDB80BC340DC07D1F000",
INIT_05 => X"FE1DFE4C080F884FE33C078F803F19F011E93ED49BE01F1A03B8972E6D20F049",
INIT_06 => X"64A08857902000DE142D4142D5030010134395D70589415002FFF800F0C38111",
INIT_07 => X"00088400092300601CE00101DE040811D919F402244293FEE00400CCB46BA4C1",
INIT_08 => X"7FA0AA08148A4000887FE0000F20C8C80D080D818FC2000000418FD08142BAD0",
INIT_09 => X"0BFA02E204D2154D28AA3FC60888D03C10415A80402847F8002458926A002E45",
INIT_0A => X"0406305587A1540231410006DFFF80540541619968C76980E914E4163D498010",
INIT_0B => X"FFFC0007C7C0140D0B50A8218102C0816040B1225C1506512C83E85500AC3A08",
INIT_0C => X"40520000141EC0000000A01000141EC0000000A01008480D3EB4A24A0C910037",
INIT_0D => X"0001A000141EC0000000A01000141EC0000000A0100100800050000000000000",
INIT_0E => X"00000000000040B000010401A0E000000000000046000002080429C000000000",
INIT_0F => X"80000340483B590000202000008402C080000000000000240801000100800060",
INIT_10 => X"28B10000001A08020002040000000020013600004414588000000D00108484C0",
INIT_11 => X"281D000000000021560002200011454000000000400902109098200000680088",
INIT_12 => X"000000008320C00000000000086016000220000120000000000082D800082000",
INIT_13 => X"D6ABC032936E43A92F2880B01F37001004B29450580000066021F6303C000408",
INIT_14 => X"45624DB481806A62840800C22800B8900042FF0180000ABFEF89250815568A8A",
INIT_15 => X"68D0068D0068D0068D0068D006A68034680300021410028450530014014002D4",
INIT_16 => X"2C989489418D13FE7F3FFD8BADB7FC4F4164A00806522C0A40A50268D0068D00",
INIT_17 => X"C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C4B1",
INIT_18 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_19 => X"2FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_1A => X"5D75D7FFEFFDF9FAF3E7E3EFFFFFFEBFD6EE7FFDF7FE78FC3CEFFDFFEA0C0060",
INIT_1B => X"EFF7FBFDFEFF7FBFDF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DD75D75D7",
INIT_1C => X"001F7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDF",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"3CF3CF75EFBD75F5FFEFFDFDF7DF7FFFFEFF9FE1F7FFBFEFDFBBFDFFD0000000",
INIT_1B => X"FE7F3F9FCFE7F3F9FCF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"0007F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"1084B030000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"6DA986092050306382C05A1C900000001FAE89016387B2A38B5000D03FA1C0C2",
INIT_05 => X"F8F92B90307F41338E303F0E07FE19C7F1FB7F289B81FB8003A396D20940C3DB",
INIT_06 => X"DF800106000FFC020004C0004C0006288004880800036002137FE3E101030222",
INIT_07 => X"000100000000000000000220000810200220620E00030BFE000181092CE7ED80",
INIT_08 => X"7E4F400000000001107E8FF90001000040100000004102200000801102448100",
INIT_09 => X"23E0FC027DF780DF74013F1C00240071E79F05888C618BA3F800599C10104903",
INIT_0A => X"040100240A808004420400202FFC3E002202021259CFDB039E00080245100000",
INIT_0B => X"FF40FFC407500020004C10060204010200810040801060C04821202001A05A00",
INIT_0C => X"00020201E04000010007400001E0400001000740000803C0616184184031010F",
INIT_0D => X"00000001E04000010007400001E04000010007400000BD0020000008001F0100",
INIT_0E => X"0200001EC00000102006E80800000010001DC0000000400D7010000008000077",
INIT_0F => X"01C200000308C50402144235400000000010003C064000C000010080BD002000",
INIT_10 => X"4000000E400000FC0010000000FC000000140403A020000007200000E8080000",
INIT_11 => X"000000001F01000014040455808000000007B00000001D010000003840000740",
INIT_12 => X"903A8000000000403C34000080001404045D00200000007C400000501001DC08",
INIT_13 => X"001A1FE004048240426200081F147FF0018C1380DA10400140640100D4080032",
INIT_14 => X"812982050800A91012494C31004124080886FE187FC301B124F2001600000000",
INIT_15 => X"1000C1000C1000C1000C1000C18006080060840477330C4889CC012188310E08",
INIT_16 => X"44602002061004A820104809402BE1900222019861D1403803800C1000C1000C",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"2FFFFFFFFFFFFFFFFF8100401004010040100401004010040100401004010040",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000100080",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"88280C4C7B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"00160090920C04800904848262220277E05152B280780D407428E723C01E1400",
INIT_05 => X"0006D46207801E400183C0707800E6000E008057641E00473C40680D32330C00",
INIT_06 => X"203F70C165000225E2C11E2C12A0D0144AC27206582C166504800000B0FC21D5",
INIT_07 => X"920CFC5E6D233B964E7CD99DFB870E1DDDD889C5FBDC440129A0604442180238",
INIT_08 => X"80B036AD23C17544C581000657A0E8E83D86F0E4A7B2D88AAAFD7FE0E1833AC5",
INIT_09 => X"C800016D82082E2081B6C0027ADA398000008A504318404005B70663212C04A0",
INIT_0A => X"4AF4AA414568729139FAD610C00001A2502440888420247041E87681008CE9AF",
INIT_0B => X"00890022B826E250B12346F1244812240912048941621804A150CA1CA45C254D",
INIT_0C => X"B2E0F1F80FA97FE0F0009E0FC40FA97FE0F0009E0FC048211E9C11C31F82E4A0",
INIT_0D => X"C3CB5F040FAB3FE0F0009E0FC40FAB3FE0F0009E0FCC42EFDFBF0AE03080E2AE",
INIT_0E => X"187806013879BA878FE807F65FBF12E0380231F0BD9E3FC08FEBD6F661C0E008",
INIT_0F => X"C83136B248831ACBFC8BBDCAB779BC699F20180309A0F83BE2B87C7C42EFDFBF",
INIT_10 => X"9947184131B59003FFEC07F00003F01FB90BE9F01FC8B38C2098DAE007F323A0",
INIT_11 => X"D065703080E29F1B2BE9F8A27E6E915C0E004C72BEC800FE7464290626D7003F",
INIT_12 => X"6F846DFC0C2352A0024B83F07F198BE9F8A0FFDA2A3C0202B8776A2FA7F023F7",
INIT_13 => X"11800014481A6105810941C5C068000CD4004C0905E52630BB1AE49C2BA7F98D",
INIT_14 => X"7E96656074EA560F0416A24844B01302A26100C4801844069B0C88881A28C141",
INIT_15 => X"E2781EA781E2781EA781E2781C33C0613C0E21020800239450116ED443C041B4",
INIT_16 => X"8112C1241140A056954AB0C280D0002020187007122C3E04E03383E2781EA781",
INIT_17 => X"1204812048120481204812048120481204812048120481204812048120481205",
INIT_18 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_19 => X"4000000000000000001204812048120481204812048120481204812048120481",
INIT_1A => X"10410411062084E57CE2641DC71C71574E09B56C74DAB16782171CF13043A85D",
INIT_1B => X"F87C3E1F0F87C3E1F04104104104104104104104104104104104104104104104",
INIT_1C => X"0007C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0",
INIT_1D => X"0000000000000000000000000187C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE500",
INIT_1E => X"BD54BAF7FFD55EF007FD75EFFFAE97555557BD75EF5D00000000000000000000",
INIT_1F => X"FFC0000AA843FE00AAFBE8B45AA803DFEFA28428B455D0017410A28428AAAA2F",
INIT_20 => X"57FFFEBAA2D5401450051401555D7FC0145F7AEBFFFF08002AA10A2AABFEAAA2",
INIT_21 => X"5D7BD755555517FFEFA280021FF082E974AA5D7BFFE000804000BAAAAAAAB455",
INIT_22 => X"A5D2EA8B45005168A10AA8028A10087FD7410557FC21555D51574AAA2FFE8B45",
INIT_23 => X"FFFFAE95410AA80000005D003FEAAFFAEBFE00A2803FEBA002A820AA0800174B",
INIT_24 => X"5EFA2AEA8A10000417410A2FFE8BEFF7FFE8B45FFFBC00005D003FF45557FC01",
INIT_25 => X"000000000000000000000000000000000000000000557DF5500003DFEFFF8417",
INIT_26 => X"12555F524AFE38B780154BAFFF1D54AF0075D75EFEBAE9554540754717F1F800",
INIT_27 => X"B6AB50B6AABDE12BEA0AF010B7D1F8F47E00A2DB45AA8A3AFD7B68E2AB78550E",
INIT_28 => X"A43FE9257F1E816D557095EAAA2D1401D500002A150038038E285D7F78FD7000",
INIT_29 => X"57545A87AAD178A8002D1D21C5E8257D5C7AA854008700249243A412EBFF5542",
INIT_2A => X"02D152A82000E3A5D2150AB8F401471EDBC0B680900AAF52B474385D75C502D1",
INIT_2B => X"D417FD7E9541242FE920AD082E10A28F6A150012A2F02AFFDF40E85F475451D5",
INIT_2C => X"55080550E87B7A405B52AAD152BD00151EAFEDB52E3F1EFFFF485A2DA3D5D24B",
INIT_2D => X"445057F40545850000000000000000000000000000000000000000000005AAF5",
INIT_2E => X"AB55F7AEAABFF5D2A81151FB8635A02FA69574BAF7D5555AF0D79D55FFA2AC97",
INIT_2F => X"34A08D46F6ABE7082AAAAF2FAC77FE00FF16565B2FA9075F4F7B3EBDF50FEAEA",
INIT_30 => X"C95256803CE3AEB038662E5D81406014D5D51F5E08A394003A908B8410E707EF",
INIT_31 => X"C0954AF0151555AF58794040077D774FAE8C798A11A0EAEF75F7AA84001A7052",
INIT_32 => X"245B4E1870108B11020AD4AA05542A0A05051023F9A9D57B63BFBF906CB45FAB",
INIT_33 => X"ABD5F5F0DA6BC9525688C1A2A0C06E9FEE5555BE48AB2A2AE0A0F20C43EAC562",
INIT_34 => X"0FF8000000FF80F55E25C00A0BA7FBED407A97F6F35F498B96BEB12DAAB77558",
INIT_35 => X"00FF8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF800000",
INIT_36 => X"000000000000000000000000000000FF8000000FF8000000FF8000000FF80000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000800000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"CA1800080848B0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000010822C00803804000001999EF9C00040B0002000001000640200001018",
INIT_05 => X"0000400244000000014200004000000004000000001000032000200002100800",
INIT_06 => X"202800208500000080412804100CB08000302220080408010000000404100844",
INIT_07 => X"25FC4C5AF6FEF002230018010860C1833C460044204C000008A0041000080008",
INIT_08 => X"0010008D22C0F55000010000524481890BC000263000188AAAA10F8C1830562B",
INIT_09 => X"041001B102002E20013600022D8819000000A000110A4000002C204000240420",
INIT_0A => X"0BE0B002605C1C1108484400C000002040040820000020104100028800002801",
INIT_0B => X"000000081001004010810510040802040102008100200800A1100707040101E2",
INIT_0C => X"10F18058000003C0F000A000C4000003C0F000A000C0000012187087010AE4B0",
INIT_0D => X"00012704000003C0F000A000C4000003C0F000A000CC4200002F08E030800000",
INIT_0E => X"1878060000000AAC00680000001F10E038000000078808C00000023461C0E000",
INIT_0F => X"4800025200040A00D000000202090C281F201803000000240218C0044200001E",
INIT_10 => X"904618400012900001EC03F000000000392100B00048230C200009A000130320",
INIT_11 => X"806070308000000961002880204A901C0E00000002C9000260640900004D0000",
INIT_12 => X"0904285C0C0312A002000000083881002880025A0A3C020000002A8400B00007",
INIT_13 => X"08400004080030008010468220A00008D0000801046004308A18500002012800",
INIT_14 => X"2200000840280206089000004090110200000000001454000200828008081110",
INIT_15 => X"A4191A4191AC191AC191A4191A00C8560C8D2910000060901010401E13405111",
INIT_16 => X"8000410410028000100800140000002004103224002006406401918C191AC191",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"0000000000000000000200802008020080200802008020080200802008020080",
INIT_1A => X"1451455901218D2C4CA2900C9249258306BABEFC54A081701C397452B4008A04",
INIT_1B => X"BADD6EB75BADD6EB755555555555555555555555555555555555555545145145",
INIT_1C => X"0005D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2EB75",
INIT_1D => X"0000000000000000000000000607FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF600",
INIT_1E => X"E80010AAAABFFFFFF803FE10F7D17FEBA55556AAAAAA80000000000000000000",
INIT_1F => X"2EBFEBAFFD555400557BD54BA5D7FFDF45A2FBD75EFA2AE97555F7FBFFF45FFA",
INIT_20 => X"A802ABEFA2D568A005D5157400AA8028AAAF7FBD54AA002A955555D7FE8ABA08",
INIT_21 => X"FFFFFDF55AAFBC0010555540010550417555AA8028BEFAAAE97555082A80000A",
INIT_22 => X"A557BD7410550428ABA5D5168ABA552EBDFEF5D7FEAA00AAAABFEAA007BC0145",
INIT_23 => X"FFFFFFEAB55557FFFEBAAAD568B45A2D5575555D7FC2155F7AEA8BEFAAAA954B",
INIT_24 => X"4AA5D7BD74000804154BA082ABFF55FFD57DF45F7D568ABAF7AABFFFF082ABFF",
INIT_25 => X"0000000000000000000000000000000000000000002EBFFEFA280021FF082E97",
INIT_26 => X"95545E175EFF57BF8FC2000BEA4BAE97F78A3FE28E3D17DEAA485FE8E02B5000",
INIT_27 => X"FD55455571E8A2A087BF8EAAEB8E0016D5D75D54BA5D7BFFF7DA2FFD55EFAAA4",
INIT_28 => X"AA07157428145A00AA8A2FBD7B6DF6AA28550E10405F7A4AFE38EAA0924921C2",
INIT_29 => X"6AAB8E971471C7010B7D168F47400A07A28415A001684104155C5B6DF6DBEFBF",
INIT_2A => X"5FD4BFBD7B6A0BF492415FC20105D24AAABF1FFBC7010FF8A38FEF557FEAB78B",
INIT_2B => X"FE38017EBA4A8EB8F6FFD5FE8B7D557495EAAA2D16D1FDBED56A55557A43DE38",
INIT_2C => X"C7AA854008700249243A417FFF41542F5D717FE2AAAA56DEBD17FE3DF7FB7FEB",
INIT_2D => X"FBA007DFCA127B8000000000000000000000000000000000000000000002A3D5",
INIT_2E => X"FFEFAAFBD55FFAA8416545A6FB60F47AF2A00010F78028B15F7823FEAAA2D57D",
INIT_2F => X"21A022A38C20B2552E975F758516AAAA0869AAAB8A7C19C55550E8574BA557BF",
INIT_30 => X"895755FFEFBCEE5FBAACB10085EE5DE10A2AEBFF55F7BAAA8565DBAC1112FFAC",
INIT_31 => X"02EABEA097BEAAFAF2863FA00DD574201E7AD1FFF5575841DE08007FC2048002",
INIT_32 => X"AF9554FF57EFBFA18D4FBFFF40FF809D4000D7FC00FC5D062BBA05ED5034472A",
INIT_33 => X"FED17DFBFF6963FCAAA2283CF14050062B0A2F7AE8B5D5D51F5E18ABD5EAFFF2",
INIT_34 => X"0000000000002CB75F7AA84001A7052C95256807DC31AA8114DE55F5BED201FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000800000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2812",
INIT_01 => X"0005A18A0849204D1CA024A542500368404000720885800802000106E4D10204",
INIT_02 => X"5C010802020408040C600850AA055254090541A111240A104A0000000908B510",
INIT_03 => X"182202210800004401060A0010041028021560A0218808002440840008C80550",
INIT_04 => X"21030A008814500120A06B0870201010258261E141A2326511024182142494D2",
INIT_05 => X"48484098142953388552102442884882B58A09291290A1120A81A3C200418DCA",
INIT_06 => X"22208802800554529001C9003A2800203120000104810100002A614008102244",
INIT_07 => X"0008040000221040408100890C0000011804480420420154000088096A0EA8C0",
INIT_08 => X"B846C0081190C105424705510A08828A0B190C0428040080A0A10F8000009200",
INIT_09 => X"20B0573165541CD54822160A89E89020AA8A80CA9D39CE215264B15818004442",
INIT_0A => X"0402100C088104010AC80005C568147007031012D40D71824114081538000048",
INIT_0B => X"550055481205100C000134128304408020C11020040244D00001306100A24600",
INIT_0C => X"00500000B01480010000A00001501480010000A0000801487334E34C1A980001",
INIT_0D => X"00012001501480010000A00000B01480010000A0000138000040000800000000",
INIT_0E => X"02000000000000A00003600180400010000000000608000A5004090008000000",
INIT_0F => X"000002400008C4000220420040800280001000000000002400000001A1000040",
INIT_10 => X"2090000000120C94000200000000000001380001C01048000000090298040440",
INIT_11 => X"2018000000000001580002508010440000000000000953008088000000481380",
INIT_12 => X"10180000820080000000000008201800024C000100000000000002E000095000",
INIT_13 => X"09130A82000C90A0000081A004342AB001720040000000000001502050000422",
INIT_14 => X"094882958000934200904407600090822085E0100D52498002B1041092001514",
INIT_15 => X"3C1011C1013C1011C10134101140801A0808AD4451394CD0391A541593C04B59",
INIT_16 => X"022810800000A0289A6D084D4021208106142034406144004041011410114101",
INIT_17 => X"4010040104411044110441100401004010040104411044110441100401004010",
INIT_18 => X"0102401024010241106411064110640102401024010441104411044110040100",
INIT_19 => X"2F81F81F83F03F03F04110641106411064010240102401024110641106411064",
INIT_1A => X"0820823047486021658010816596597700138D70C030B542923650C7D0002281",
INIT_1B => X"944A25128944A251282082082082082082082082082082082082082082082082",
INIT_1C => X"F804A25128944A25128944A25128944A25128944A25128944A25128944A25128",
INIT_1D => X"0000000000000000000000000787C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF871",
INIT_1E => X"5420AAAA843DFFFAAD1554005D7FD74AA0004001550000000000000000000000",
INIT_1F => X"2EBFF45AAAAA8A10A2AE80010A2AA975FF5D003FE10F7D17FEBAF7D5420AA085",
INIT_20 => X"D7FFFF45A2AA975EFA2FFD7555FFFBFFF45AAFBC20AAF7D1575EF55517DF555D",
INIT_21 => X"AAAE95555552E974105D517DF55AAAAAABEFAAD1575EFAAAE974AA5D51554BA5",
INIT_22 => X"F552E82010F7AABFE10FFD542145FFD5554AA555555555557FE8ABA082EBFFFF",
INIT_23 => X"EFF7FBC0010AA802ABEFAAD540000FFD540000AA802AABAF7FFC2010AAAE821E",
INIT_24 => X"555AA8028BEFAAAE821550851420AA002E800AA08042AB45007FC00BAFFD168B",
INIT_25 => X"0000000000000000000000000000000000000000002E80010555540010550417",
INIT_26 => X"7DEAAE95F40002157F470AABE803AE97A2DF55400557FD54AA1D04001C515000",
INIT_27 => X"E105EF55517DFC5552ABDF45B6AEAFFD5F7A482000BEAE905C755003FE28E3D1",
INIT_28 => X"A4070BA5FD0154BA5D7BFAF7DA2AE955EFAAA495545E3F5EFF57F7FE80082FFD",
INIT_29 => X"571E8AAF082AB8EAAEB8E0016D5D2A924105D5B7FF7DB6AAAABC7BEDB505EFBE",
INIT_2A => X"E80495038AAAEAF1D7410E80000FF8438E00B6DF68FEF4871D24BA495B5556D5",
INIT_2B => X"80071ED1EFEAF1EFFFDEAD1C5010AA8E2FBD7B6DF47A00EBDB50000A380AAE28",
INIT_2C => X"28415A001684104155C5B68E2DBEFBFFBC703AE2DF42AAA002A851C214003FF6",
INIT_2D => X"4AA550002155510000000000000000000000000000000000000000000002087A",
INIT_2E => X"215555003FEAAAAD57DEBAA2FDDC01051FBD74BAF7802AB05AAFBD5400557BD5",
INIT_2F => X"60F47AF7FC20B2F7FBC015D58517FF555D2ABDF55F782BEB47AFAD00010F7AA8",
INIT_30 => X"22A955FFFFC20FFF3AE544108410174BA557BEABEFAAEBD55FFAA1456547A2D3",
INIT_31 => X"D4420BA547FD75FF58516AAAA0828AAAB4A78016545540400010557BFDFFFF78",
INIT_32 => X"FFBD550AAFACAAA122AA8954BAA2AE9D545002A800A8FF862BA00F2F9E8F0050",
INIT_33 => X"002E954505C417FFFF08555555BAAD335B57AB5155400A2AEBFF45FFFB404007",
INIT_34 => X"000000000000061DE08007FC2048002895755FFAEBCFE57BBA57002DF3C4AAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000001000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B815602110494074133520400E02B92206",
INIT_01 => X"014C9BC048800168240442C99E004B61404040028804A0080A000516A0990A08",
INIT_02 => X"4809A900031800444440589866E331352180D468B8000E600C0081110B802CD0",
INIT_03 => X"DA16C0200C0001423583480408D60520320066810A80881068A808029C856330",
INIT_04 => X"2088681DA82740EC92307364B37569100A84E1E11C251210990040420E005A48",
INIT_05 => X"2D284A102414411A314A0A02C18C01B9854368280A506902018C2442484038D1",
INIT_06 => X"23600016801CCCAA9061C9061C0D0080001005210C8761001166CCC40C110826",
INIT_07 => X"0178045800B6540063000889082040A13A0716042440833280038C89904E6400",
INIT_08 => X"D20A480810804451421D1CC8024481994B5500061000088000A10F840854973A",
INIT_09 => X"2079CCB035E03CCC5D2A35620988100A698761C0953B6E84C82C404018304D42",
INIT_0A => X"070070202A90340440C80004CCE4CC1042061913208CE8024380880820010040",
INIT_0B => X"3302CCC01300104018900402870C4287214210E114200410EC20242D01015E84",
INIT_0C => X"4801000180148000000800100040148000000800100401C33249049051218073",
INIT_0D => X"04008001001480000008001000E014800000080010001C000040000000000000",
INIT_0E => X"0000000000004408000068018040000000000001400800091004090000000000",
INIT_0F => X"00004100812644000004400140800280000000000002000008008000B0000040",
INIT_10 => X"20900000020800CC0002000000000020400800030010480000010400C8040440",
INIT_11 => X"2018000000000060080004418010440000000000410015008088000008200540",
INIT_12 => X"80188000820080000000000100400800041C0001000000000000902000014C00",
INIT_13 => X"284B264208448260E27285A23224E660084208410000004444000E0000000020",
INIT_14 => X"0840024D810283021280400720C0348002854C001CC3158026A2040028090441",
INIT_15 => X"80901A0901A09018090188901A248054480C0C0041116DD0115E011599641E59",
INIT_16 => X"C6C8408514028028D06C0C5D20030BA1010021B000020402400501A090180901",
INIT_17 => X"4290C4290843908439084390843908439084390C4290C4290C4290C4290C4690",
INIT_18 => X"290C4210E4290C4310A439084310A439084310A4390C4290C4290C4290C4290C",
INIT_19 => X"5D54AAB556AA9556AAC310A439084310A439084310A439084210E4290C4210E4",
INIT_1A => X"0820825103A1600054C0F4012492490300C78C706428A1411133586294020A90",
INIT_1B => X"D4EA753A9D4EA753A92492492492492492492492492492492492492482082082",
INIT_1C => X"8086A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A353A9",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE024",
INIT_1E => X"5421EFAAFFD54AAF7D168B45AAAABDF5500002AA100000000000000000000000",
INIT_1F => X"043DF45FFD168AAA0855420AAAA843DFFFAAD1554005D7FD74AAA28400155005",
INIT_20 => X"2AA955FF5D003FE10F7803FEBAFFD5420AA080400155AAD5554AAF7802AB4500",
INIT_21 => X"AA8028B45A2AE82155A2FBFFEBA0800021550855555FFAA84001FFAAAE80010A",
INIT_22 => X"0085168ABAFFFBD54BAAAAE97400A2FBC20AAA284175EF55517DF555D2EBFE00",
INIT_23 => X"55AAAA954AA5D7FFFF45AAAA975EF007BD7555FFFBFDF55AAFBD55EF5D2EBFE1",
INIT_24 => X"BEFAAD1575EFAAAE974AA5D00175555D0015410F7AAAAAAA55043DE00FFFFD55",
INIT_25 => X"00000000000000000000000000000000000000000004174105D517DF55AAAAAA",
INIT_26 => X"D54AABC04001C51551471D7AAF1D05D2EBD56DB7DBEAEBFF551C042AA101D000",
INIT_27 => X"B50492EB842FB5508043FF55EBD56ABD75D5B470AABE8A3AFD7A2DF55400557F",
INIT_28 => X"8E82557FD2082000BEAE905C755003FE28E3D17DEAAEBDF40002550F47155AAD",
INIT_29 => X"5517DF40552ABDF45B6AEAFFD5F7A48017DAAFFFAE821C0A0717D1C5B575FFB6",
INIT_2A => X"F7D5C55D7492E90E3808756DA92EBFFD74BAE3AE85480FFFFC00AABE8E105C75",
INIT_2B => X"241043AE10EAF5C5547FF80954AA5D7FFAF7DA2AE905EF0075D5545E3F5EFF57",
INIT_2C => X"105D5B7FF7DB6AAAABC7BEDB505EFBEF5C7092FF801756D490A10438EBA4B8E9",
INIT_2D => X"F555D0028A00510000000000000000000000000000000000000000000000E124",
INIT_2E => X"8B45AAFBD54005D7BD54AAF78002155515157555AAD142040A2D57FFFFFFAEBF",
INIT_2F => X"DC01051AE955F7AAFBC0000AF843FF5500003FF55AAFD6AB455157D74BAF7AAA",
INIT_30 => X"E955FF557BD74EFFBACD41577B8400010F7AA8215555003FEAAAAC53DEB8A2FD",
INIT_31 => X"FEC20BAF7AA8015558517FF555D2ABDF51F782BCB47ABAE801FFAAFBEAA105D2",
INIT_32 => X"8554214FA2D3EAF57AFFDD7555082AA0AAA00557FEA8A2FDD64BAAF8282012AF",
INIT_33 => X"082A820AAAB842AA00000028AB0AAFF48547AE04174BA557BEABEFA2AA951FF8",
INIT_34 => X"0000000000002A80010557BFDFFFF7822A955FFFFC21FFF3BE40412DE02955FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000800000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303000048B3532C82D04A16002",
INIT_01 => X"210399800808004C1C20650E1E104368403008418984014902030006A8910200",
INIT_02 => X"480108A200000000444148E41E80F00A4104311868200200080000000988A390",
INIT_03 => X"0CA08220080000D004260A0240109028270012603000000030808C4208C000F0",
INIT_04 => X"4403A609A055306BC2C0735810CEE5100A0A48E16B8370E3808241D03845D002",
INIT_05 => X"ECE8698800791403AD3038AE079059A790E245A19A41E4120BAB86C00001D312",
INIT_06 => X"23208806000C3D220023C0021A21008891048C00040341121661E3C10000A064",
INIT_07 => X"0008045000220440000000090800102118400204A04100F040018019004B8001",
INIT_08 => X"0E11400810906441123323C0424190880B0108002000000880810F9002041200",
INIT_09 => X"22003C2309671584786E0F5A88889031EF9F05D884794FA03A24781810106D02",
INIT_0A => X"0409400E4282A00142400004DC3C82400702003200872003FB14080828400010",
INIT_0B => X"F050C3C00095000C008135040002010100800040001400C00401208800F01A14",
INIT_0C => X"08000002E0100000000800000220100000000800000001C87261C51C42390240",
INIT_0D => X"0400000280100000000800000360100000000800000035100040000000000000",
INIT_0E => X"00000000000004000000D8008000000000000001000000155000080000000000",
INIT_0F => X"000040000120EC00004002214000008000000000000200000000000094100040",
INIT_10 => X"001000000200050C000200000000000040080005800008000001000168000040",
INIT_11 => X"000800000000004008000448000040000000000001003C000008000008000D00",
INIT_12 => X"800800000000800000000001000008000017000100000000000010200002C800",
INIT_13 => X"150F5E0400101000227200800E271E00288400800208004C04C0080000000052",
INIT_14 => X"818082450000920280C544310041B408880EC51060461589225100063E9012D6",
INIT_15 => X"1410C3410C1410C1410C3410C100869A08618C00772201D899BA003591510A59",
INIT_16 => X"44E0110004480020986D4815044369A00006203041C3443043010C5410C3410C",
INIT_17 => X"0080001002008040100200800000060180000006008000100600804000020180",
INIT_18 => X"0000010060080201800000040100201802008040100201804000020180001006",
INIT_19 => X"64B261934D964C32698080401000000060080601800000040000201806008000",
INIT_1A => X"1451457A604C8D0C28A280CD145144C1863807E0500014385DAF345041488280",
INIT_1B => X"1A8D46A351A8D46A355555555555555555555555555555555555555545145145",
INIT_1C => X"1F60D068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D06A35",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE077",
INIT_1E => X"02ABFF087FFDF5508003FEBA087FD54BAAA84154005500000000000000000000",
INIT_1F => X"2EBFF5500003DF455555421EFAAFFD54AAF7D168B45AAAABDF55A2802AA10000",
INIT_20 => X"A843DFFFAAD1554005D7FD74AAAA840015500002AABA082E954005500021FF5D",
INIT_21 => X"FFD168BEF080028BFF0855555455500174BAA2AABDE0055517FF555555420AAA",
INIT_22 => X"0085168ABA0055574BA5555554BA5D0400155AAD1554AAF7802AB4500043DF45",
INIT_23 => X"AA5D0400010A2AA955FF55003FE10F7803FEBAFFD5420BA085168A00007BFDE1",
INIT_24 => X"1550855555FFAA84001FFAAFBEAB45002A97545F7D1555EF55043DF5555517DE",
INIT_25 => X"0000000000000000000000000000000000000000002A82155A2FBFFEBA080002",
INIT_26 => X"BFF55BC042AA101D0A28BC7007FFDF45080A3AEAA007BD2482BE84124285C000",
INIT_27 => X"4974004100021FF492AB8F7D1C0438E381451471D7AAFBD0492EBD56DB7DBEAE",
INIT_28 => X"557AFED1C5F470AABE8A3AFD7A2DF55400557FD54AABE84001C5550A28ABA142",
INIT_29 => X"B842FB5508043FF55EBD56ABD75D0428BEF005557545490012482B6A0BAE2849",
INIT_2A => X"557F6DA101475FDE10145F68A921C55504924955524AA140E0717DAADB50492E",
INIT_2B => X"F5D043AF6D405F78E3A1C2002000BEAA905C755003FE28E3803DEAAEBDF40002",
INIT_2C => X"7DAAFFFAE821C0A0717D1C5B575FFB6DF425575D7BEFB55002097555FFD5401E",
INIT_2D => X"010F784000AA5900000000000000000000000000000000000000000000020801",
INIT_2E => X"2000A2D57FFFFF7AEBFF55FF8028A00512EAAB45007FFFF55082EA8AAA087FC2",
INIT_2F => X"02155512AAAA085D04174100800021FF002EA8BEF5D0428ABA595557555AAFBC",
INIT_30 => X"402000FF802ABAA04552ABFF597FD74BAF7AAA8B45AAFBD54005D7BD54AAF780",
INIT_31 => X"2F955FFAAFBC0000AF843FF5500003FF55AAFD6AB4551002ABEF005555555000",
INIT_32 => X"A843DEB0A2FD5600051537DE005D557DE005D7BE8AA85555400100879560AA59",
INIT_33 => X"000417545FFD5421FF5D0428BEF0079FCABA598400010F7AA8215555003FEAAA",
INIT_34 => X"00000000000004001FFAAFBEAA105D2E955FF557BD75EFFBBCD415521FBFDF45",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000001000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB0A0791B1B41694368283C81F9996A091A32152007AB37B20E07C0C1E002",
INIT_01 => X"881FBC449030884C446A00000034824841280A00084000C8C212812EEA953231",
INIT_02 => X"C809AD5CB118E640A4F408FC011FF0002080000082CCC66609DB7DDDCB1F2036",
INIT_03 => X"4A100E4D3E4C90D290831C824A4204720B20048A88800000B8E0F91028C5500E",
INIT_04 => X"00144884922644001914830051110A71E03040F0105B001C662AE22DC08A3408",
INIT_05 => X"120340220B88820041CDC451B860A6506BEBD08265AE105714505F0152122449",
INIT_06 => X"207F7890752C037372A1D72A398CD084C890EA2950A37E270660182C0D2C8080",
INIT_07 => X"9378355E64B66F96231CC81D2DAB468D38C601C5FFF54FF1C9A46490261C4B39",
INIT_08 => X"7F105CAD1089654115814FC60284A1A93B46F4621030C800001D7FA56891162E",
INIT_09 => X"E00A003C832D25328526C082DF9AB88C104024C09639441807B78661090C24A1",
INIT_0A => X"4FD32A2E2A9992944AF2D611C3FC01B2152109204C28B67061EC928920C569E7",
INIT_0B => X"F0313FE92C22F21CA0B363C0A242502028901408154218144D712664A5F15AC1",
INIT_0C => X"B2F0F1E01BE53FE1F000BE0FC41BE53FE1F000BE0FC80020130841840308653F",
INIT_0D => X"C3CB7F041BE1BFE1F000BE0FC41BE1BFE1F000BE0FCD806FFFAF0AE83080E2AE",
INIT_0E => X"1A7806013879BAA78FC103FF5F1F12F0380231F0BF9E3F02A7FFD63669C0E008",
INIT_0F => X"483136F200A822CBACAB9DDEB7F9BC291F30180309A0F83FE2B87C7D006FFF9F",
INIT_10 => X"D1C6184131B7980DFFFC03F00003F01FB931E9C1DBF8A30C2098DBE2FF7F2320",
INIT_11 => X"F060703080E29F1B71E9F6427EFE901C0E004C72BEC95FEF64E4090626DF15B7",
INIT_12 => X"EFAC6DFC8C0312A0024B83F07F3991E9F21DFFFA0A3C0202B8776AC7A7C9CBFF",
INIT_13 => X"88F4C1C64044A264601144C5F1787E1C812A510885C56620590350ACD3A7D5B7",
INIT_14 => X"9054204DF56A974F92C3E20F24301300082C38C4184F10281204888298284616",
INIT_15 => X"A238CE238C8238CE238CA238CC11C6411C670C10EB4124C2B3923BF5C9710C59",
INIT_16 => X"276A11A03444922898494C5504008401230E71B3100C1634E3138C8238CC238C",
INIT_17 => X"5094650142511405194450942511425114450944519425114250144519405194",
INIT_18 => X"0944509465114251146501465014051944509445094051942501465014051940",
INIT_19 => X"2124B2DA6924965B4D5094450940519425014650142511425014450944519405",
INIT_1A => X"7DF7DF6FEFFCFDFD796ED1DCF3CF3DF6CE7F7B9DB7FF3A7E1FBC6DB7E8418A88",
INIT_1B => X"EEF77BBDDEEF77BBDDF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF",
INIT_1C => X"024F77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDD",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE056",
INIT_1E => X"5574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF80000000000000000000",
INIT_1F => X"D16AABAF7AAA8BFFAA802ABFF087FFDF5508003FEBA087FD54BA080415400555",
INIT_20 => X"AFFD54AAF7D168B45AAAABDF55AA802AA1000003FEBA00002AABA5D2EBFEBAAA",
INIT_21 => X"00003DE005555575EFA2D142145A2FFE8B45FF80001555D2E955FFFFD5421EFA",
INIT_22 => X"F5D7FC00BA5D5568AAAF7AAAAAAAAA802AABA082E954005500021FF5D2EBFF55",
INIT_23 => X"BAFFD5420AAAA843DFFFAAD1554005D7FD74AAAA840014500517FFEF007BEABF",
INIT_24 => X"4BAA2AABDE0055517FF555504154BAA2FBEAA105D2E97410FFD16AAAA5D2ABDE",
INIT_25 => X"0000000000000000000000000000000000000000000028BFF085555545550017",
INIT_26 => X"D24821E84124285C51574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7800",
INIT_27 => X"428A925D2AB8EBABEDB6AA92F7AAA8BC7B68A28BC70075FDF45080A3AEAA007B",
INIT_28 => X"2A925FFFFD1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0A38EBA1C0",
INIT_29 => X"100021FF492AB8F7D1C0438E38145B575EFA2DB45145B6F5EFB6DF78E0514555",
INIT_2A => X"55517DFC70875EABC7557FC20AA415F68AAAF7AAAAA82BE8A28A921424974004",
INIT_2B => X"0FFDB6FABA542ABAE2AF7DF470AABE8A3AFD7A2DF55400557FD54AABE84001C5",
INIT_2C => X"EF005557545490012482B6A0BAE2849043AFED1C0E10492B6FFEFA105D2A9541",
INIT_2D => X"E005D2AAABEFFB8000000000000000000000000000000000000000000000428B",
INIT_2E => X"FF55082EA8AAA087FC20105504000AA5955554BAFFAEBDE10F7FBFDEBA007BFD",
INIT_2F => X"28A00512AA8AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3AAAAB4500557",
INIT_30 => X"57FFEFFFAA97545552A821EFFBD557555AAFBC2000A2D57FFFFF7AEBFF55FF80",
INIT_31 => X"AAAAA005D04174100800021FF002EA8BEF5D0428ABA597FD55FFA2FFD5555FFD",
INIT_32 => X"D7BD54AAF7800015551517DF45005168B55557FC0012087FEAABAF7AAAAA10F3",
INIT_33 => X"FFFFFFE005D2A95410F7FFFFEBA5D2EA8ABAFBFFD74BAF7AAA8B45AAFBD54005",
INIT_34 => X"000000000000002ABEF005555555000402000FF802AAAA04452ABFF592E80010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000006000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C030028180004003220200403302301C0381A0082",
INIT_01 => X"A74041C838394848188160000C42426041000000090800090210000008510200",
INIT_02 => X"080108200C1000004465580000C0080100000000010432400800800009882050",
INIT_03 => X"080200010C234040842248600210812183806584488000103080014E88C10000",
INIT_04 => X"0040584288A6C210003120000000001002A0E8A910A072101000400A00203040",
INIT_05 => X"04096A019400C118414A00014000002014100128005004020010A0C044C02800",
INIT_06 => X"20200A301223FC029931E9931900002224240249A6D3E808D51FE00909108222",
INIT_07 => X"0008040000220001820000010C0810211A440014A040200E8240089000080002",
INIT_08 => X"0040081A08944010007FA038020080880B0104182000000000090F8102041320",
INIT_09 => X"17E2FD200240B4A409223F020888100808200450001A401BF82C21185C81744A",
INIT_0A => X"0602A0244285180542402180D001BE1907939120000020044184890800011000",
INIT_0B => X"0F0400091081190E4490A502D2A36951B428DB14A688051A5E21214601A01A22",
INIT_0C => X"455D0018101480000000A01034101480000000A01033A0081300000000001880",
INIT_0D => X"0001A0F4101480000000A01034101480000000A0103142000040000000000000",
INIT_0E => X"00000000000041E8002900018040000000000000466800C20004090000000000",
INIT_0F => X"0000034D242C2000502000000080028000000000000000240946800142000040",
INIT_10 => X"20900000001A60F0000200000000002007F000322010480000000D1A00040440",
INIT_11 => X"2018000000000025D00008958010440000000000403F4000808800000068D240",
INIT_12 => X"101280008200800000000000086670000CC0000100000000000087C000301400",
INIT_13 => X"C8B5800720849A72700094A2202301F05103202420000810C219500150002800",
INIT_14 => X"81088A454110030212C140813204D0A0888C000118471DE126805432A62A1586",
INIT_15 => X"4096C4096C2096C2096C6096C444B6004B600C446B0104D09190013589701C11",
INIT_16 => X"108D19D1804A8000904C421852240821978221B0044245B25B456C0096C0096C",
INIT_17 => X"69DA368DA1695A568DA3685A1695A768DA3685A569DA768DA1685A569DA76C5A",
INIT_18 => X"85A569DA1685A369DA5695A368DA169DA7695A168DA3695A5695A368DA3695A5",
INIT_19 => X"7638C31C71C718638E685A569DA7685A368DA5695A768DA1685A7695A168DA36",
INIT_1A => X"1C71C73B676CEDED7DE2F4DDF7DF7DF7CE7F8FF0F4FA957FCF9F7CF7F40A0010",
INIT_1B => X"FE7F3F9FCFE7F3F9FC71C71C71C71C71C71C71C71C71C71C71C71C71C71C71C7",
INIT_1C => X"2BE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"0000000000000000000000000607C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF019",
INIT_1E => X"43DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFF80000000000000000000",
INIT_1F => X"D17DEBA0855421455555574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF8",
INIT_20 => X"87FFDF5508003FEBA087FD54BA000415400550428AAAAA84021FF007BD54BAAA",
INIT_21 => X"F7AAA8BFFAAD1554BA002A95555A28417400AAFBE8ABAF7FFD54AAAA802ABFF0",
INIT_22 => X"0FFFBD5545080417555A2D17FE1000003FEBA00002AABA5D2EBFEBAAAD16AABA",
INIT_23 => X"FFFFD5421EFAAFFD54AAF7D168B45AAAABDF55AA802AA100000001EF087FEAA0",
INIT_24 => X"B45FF80001555D2E955FFFF843DEAAA2803DFEF0855401FF082EA8B555D7FC21",
INIT_25 => X"00000000000000000000000000000000000000000055575EFA2D142145A2FFE8",
INIT_26 => X"6FA92552AB8FEFF78E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FF800",
INIT_27 => X"E001EF147BD2482BED57AE921451421555551574BAB68A2DA00FFFFFFE38085F",
INIT_28 => X"FFD24BAB68A28BC70075FDF45080A3AEAA007BD24821C04124281C0E2DA82BE8",
INIT_29 => X"D2AB8EBABEDB6AA92F7AAA8BC7B6D5524AA14209557DA28E15400BEF1EFA92FF",
INIT_2A => X"5D0E071FF0071EDA38F7F1D5555000417545B6D178E281C0A38EBA1C0428A925",
INIT_2B => X"70824A8B555C7FC2147F7D1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA10",
INIT_2C => X"EFA2DB45145B6F5EFB6DF78E05145552A925FFFF8E3DE82BE8E38FFF0851401C",
INIT_2D => X"000557FE8A00F38000000000000000000000000000000000000000000005B575",
INIT_2E => X"DE10F7FBFDEBA007BFDE005D2AAABEFFBAABDFEFAAFBC00BA007BC0000FFD542",
INIT_2F => X"000AA592ABFE00F7AA821FF557FC0010F7D168A105D55421455155554BAFFAEB",
INIT_30 => X"E95410F7D57DE00FFFBC00AAFBAAAAB4500557FF55082EA8AAA087FC20105504",
INIT_31 => X"2AA8AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3D5400BA5504155EFAAA",
INIT_32 => X"7AEBFF55FF8028A00512E975FF08557FEAAF7D157545080417545F7D56AAAA59",
INIT_33 => X"F7AAAABEF005542155000028B555D7FC2145F3D557555AAFBC2000A2D57FFFFF",
INIT_34 => X"0000000000007FD55FFA2FFD5555FFD57FFEFFFAA97545552A821EFFBAABDE00",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000004800000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992006",
INIT_01 => X"A34009C0383848481C00E0000E01426040000000080000080200010000510204",
INIT_02 => X"4801082048100000446558000080000041000000000622400800000009000010",
INIT_03 => X"080001038CA14840842248400210812102000400088000003080014688800000",
INIT_04 => X"000040048106000040120000000000100220C8A5108032140004500800603000",
INIT_05 => X"04096A009000410041480081000000201000012800400022801080C0C0C82000",
INIT_06 => X"232086381A8001220021E0021803002224240248040360889100100909000222",
INIT_07 => X"0008055000220409020000090C0810211A04001420602000D2500810000C4903",
INIT_08 => X"8040491A809041100001400042409098090006102000000000010F8102041320",
INIT_09 => X"340C013102002420012200820D89140800004010900A4010002C8118D0024412",
INIT_0A => X"A221A5000800914000400888C00100200B0310200008B2066313894800631400",
INIT_0B => X"0010000800010004088105020100008000400120800000200404002450004000",
INIT_0C => X"4409081C1000000000F001F02C1000000000F001F021141A12000000000010B0",
INIT_0D => X"383480CC1000000000F001F02C1000000000F001F023420000000004C3201C51",
INIT_0E => X"00019860078641084039000000000002C0E00E0E404900E200000000000B0380",
INIT_0F => X"120C8908146000105120000000000004004160C0301D07001D04820342000000",
INIT_10 => X"000021908C4842FC000000030F000FE00600103BA0000010C8462414E8000006",
INIT_11 => X"000004C3201C60A400100DD5800000013098038D40309D000000C2419120A740",
INIT_12 => X"901A800030040902C0807C0E00C440100DDD000000411C81078884004035DC00",
INIT_13 => X"140A000410401400201020820022000250400040002211148019064200402A32",
INIT_14 => X"01889A4543148282A01415B04009904A80890033679459A926801054001C0050",
INIT_15 => X"159201592055920559205592070C901AC901A100804000801210541403C05130",
INIT_16 => X"2460010004428008904C085D44200D8001112804CDE1C483480D201592015920",
INIT_17 => X"0080200806008020000000004000020080200802000000000000000008020480",
INIT_18 => X"1000008020080000000000020080200000000000080600802008000000400000",
INIT_19 => X"5841040002082080000180200000000020180200800000000100200802000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000005428A94",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"E480000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE031",
INIT_1E => X"BC00AAF7D5575455D557DFEF002AAAB55002E820AAAA80000000000000000000",
INIT_1F => X"AEAAB55007FD74AAAA843DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFF",
INIT_20 => X"2802AA10FFFFFDE0008556AABA5D2ABFFEFFFAAAAAAAF7D57FFEFF7D555555A2",
INIT_21 => X"085542145552ABDFEFFFAA801EFFFFBFDF550000175555504175450055574AAA",
INIT_22 => X"0082A975EF00003DF55555168A00000428AAAAA84021FF007BD54BAAAD17DEBA",
INIT_23 => X"AAFF802ABFF087FFDF5508003FEBA087FD54BA000415400557BD74BAFFD14000",
INIT_24 => X"400AAFBE8ABAF7FFD54AAAAAEA8ABA55557FEAAA2843FF55A2AEA8B55AAAABDE",
INIT_25 => X"00000000000000000000000000000000000000000051554BA002A95555A28417",
INIT_26 => X"C20825D7FE8A92FFFFC70BAE3D155555415178FD7082EAAB550820870BAAA800",
INIT_27 => X"578FFFEBD55557DBEA4AFB550871D7482AA8E3DFFFAAFFD04AA415B52492B6F5",
INIT_28 => X"0E175550051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7A0ADABAEBD",
INIT_29 => X"47BD2482BED57AE921451421555524BDFD7FFA4801D7F7F5FDF55000E1754541",
INIT_2A => X"1C7BD2482E3D1450381C20905EF08003AF55415F6DA38080E2DA82BE8E001EF1",
INIT_2B => X"5BEAAAFB55ABA0BDE02EB8A28BC70075FDF45080A3AEAA007BD24821C0412428",
INIT_2C => X"AA14209557DA28E15400BEF1EFA92FFFFD24BAB6A4A8A82495F78E92AA843DF4",
INIT_2D => X"B450800174BAA680000000000000000000000000000000000000000000055524",
INIT_2E => X"00BA007BC0000FFD542000557FE8A00F3FFD54BAAAD15754508556AB45002AA8",
INIT_2F => X"AABEFFB803DEAAAAD56ABEFAAD5575EFF7803DF45085557410AEAABDFEFAAFBC",
INIT_30 => X"57FF55082E97555002E955550C55554BAFFAEBDE10F7FBFDEBA007BFDE005D2A",
INIT_31 => X"2ABFE00F7AA821FF557FC0010F7D168A105D554214551003FF45FF8400145FFD",
INIT_32 => X"87FC20105504000AA597FC2010A2D1554AA5500021EF000028B55087BFDEBA04",
INIT_33 => X"007FE8A00A2803FF45F7AABDF55AA843FE10AEAAAAB4500557FF55082EA8AAA0",
INIT_34 => X"00000000000055400BA5504155EFAAAE95410F7D57DE00FFFBC00AAFB8028A00",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"A140084000080048040100000202026040000000180800080200010048510204",
INIT_02 => X"080108000090000004655C000080000051000000000402400800000009000010",
INIT_03 => X"0000000100300C40842240000210810002800584488000103080894288800000",
INIT_04 => X"0002584280A2C21000110300100000100220C8C910A032541000090A00643000",
INIT_05 => X"04092A001400D100410A002140004020140001A9005000004810A1C0044D2800",
INIT_06 => X"0360000010EFFD229911C9911820002080258A09A2D3E102137FE0094910A222",
INIT_07 => X"0000004000220400120000090C0810210A040034A040000046180810000C4907",
INIT_08 => X"80404050D88C24510001400042008088090004012000000000010F8102041320",
INIT_09 => X"20080120024030A4090200828C880208002044C0843B44100228A1585C81740A",
INIT_0A => X"142180860A84802042C82180D0010039039390200008B20E2300086800400640",
INIT_0B => X"003000091084190644810502D0A16850B4285B14A688011A1409212008F05E20",
INIT_0C => X"400104080010001E0FF00010000010001E0FF0001002200A1300000000000080",
INIT_0D => X"000080000010001E0FF00010000010001E0FF000100440000040F517CF600000",
INIT_0E => X"E587F9E000004008100800008000ED0FC7E000004000804000000809963F1F80",
INIT_0F => X"36000100202C0020100000000802419660CFE7C0F00000000800810040000040",
INIT_10 => X"0618E7B0000800000003F80FFF0000200018021000030C73D80004000000585F",
INIT_11 => X"078A8FCF600000201802008001006AA3F1F80000400000000B0BD6C000200000",
INIT_12 => X"0041120370DCAD1FC18000000040180200800005D5C3FD800000806008100000",
INIT_13 => X"48A480072284983230101402200200111103202420000880C218000150100800",
INIT_14 => X"2B888A4500048240C08400843204502000890001000415E12480003002944281",
INIT_15 => X"0480004800048000480004800004002240020854884000901212140011C01079",
INIT_16 => X"346D19D1A4C08028904C4E1D7224086590800420044040020004004480004800",
INIT_17 => X"68DA368DA368DA368DA368DA368DA1685A1685A1685A1685A1685A168DA36CDA",
INIT_18 => X"8DA3685A1685A1685A1685A368DA368DA368DA3685A1685A1685A1685A1685A1",
INIT_19 => X"40000000000000000068DA368DA368DA1685A1685A1685A1685A368DA368DA36",
INIT_1A => X"3CF3CF6FE23CCD8D00A281F5B2DB2CA78A543EBC57A10A245DA975D640088884",
INIT_1B => X"3E1F0F87C3E1F0F87CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"5DA9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0F87C",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00B",
INIT_1E => X"40000000043DF55087BC01EF007FD75FFFF84000AAFF80000000000000000000",
INIT_1F => X"2EBFE10A28028AAAAAFBC00AAF7D5575455D557DFEF002AAAB55002E820AAAA8",
INIT_20 => X"2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFAA95545552ABFE00087BC00AA08",
INIT_21 => X"007FD74AAAAD57FF45002A975FF007BE8BFFA2FBFFFFFAAD5400AAFF843DFEFA",
INIT_22 => X"5AAFBE8A00082A97410F7D5555EFAAAAAAAAAF7D57FFEFF7D555555A2AEAAB55",
INIT_23 => X"450055574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFFAA8200055555554",
INIT_24 => X"F55000017555550417545000015545087BC2010AAD54014500516ABFFA2AABDF",
INIT_25 => X"0000000000000000000000000000000000000000002ABDFEFFFAA801EFFFFBFD",
INIT_26 => X"AAB550820870BAAA8407000140038F450075C71FF087BD75D7FF84050BAEB800",
INIT_27 => X"AB8E10007FC50BA002ABFE00AA8A2AABABEFFC70BAE3D155555415178FD7082E",
INIT_28 => X"DB45082EB8E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFA497545552",
INIT_29 => X"BD55557DBEA4AFB550871D7482AAD17DF451C24955EF0875EFBD7B6F1FFFC7BE",
INIT_2A => X"F7AA87000415B5057DAAFBE8A10082092410EBD5505EFB6A0ADABAEBD578FFFE",
INIT_2B => X"D005B6ABC7B6AABFFED0051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEF",
INIT_2C => X"D7FFA4801D7F7F5FDF55000E17545410E17555000E17545007BC0000BED14217",
INIT_2D => X"555F784174AAA280000000000000000000000000000000000000000000024BDF",
INIT_2E => X"754508556AB45002AA8B450800174BAA684174105D042AB550055555FF007BD7",
INIT_2F => X"E8A00F384175555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7FFD54BAAAD15",
INIT_30 => X"57DF55FFD57DF55FFFBD5400A2AABDFEFAAFBC00BA007BC0000FFD542000557F",
INIT_31 => X"803DEAAAAD56ABEFAAD5575EFF7803DF45085557410AED17FF455D04155FF005",
INIT_32 => X"07BFDE005D2AAABEFFBAE97410087BC21EFA2FFEAA00000002010A2D5421FFFF",
INIT_33 => X"087BC0010FFD1401EF087FE8B55FFAEBDFEF0855554BAFFAEBDE10F7FBFDEBA0",
INIT_34 => X"000000000000003FF45FF8400145FFD57FF55082E97555002E955550C2E95555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000002000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000006",
INIT_01 => X"0000098218302849180060000C004260413C0A61590001D90213C80000110200",
INIT_02 => X"680108220010000054400C00008000004100000001200240080080000908A011",
INIT_03 => X"000A0000040020400002021000000008428065044880001030818C0008C10000",
INIT_04 => X"00005042882A8210003000000800001000806080100040140080040800003140",
INIT_05 => X"0400000840000098410800010001002000000000004000002010000040002000",
INIT_06 => X"03600810100001220911E0911902000020200200A253E8000C0010080800004C",
INIT_07 => X"000408C0002204400200000B080000010C040004A0400000C0000810000C5901",
INIT_08 => X"000008002A84300000014000C2008088090008002000000000030F8000001220",
INIT_09 => X"0008012100000200001200820888010800200000000840100028800004801440",
INIT_0A => X"000090220000040400480000D0010009049090200008B2022384800802010000",
INIT_0B => X"001000090001090A4C81240050A328519428CA14328C840A5820000101500400",
INIT_0C => X"00510008100400000000A00000100400000000A00000000A12000000000000B0",
INIT_0D => X"00012000100080000000A00000100080000000A0000540000000000000000000",
INIT_0E => X"00000000000000A8000900010000000000000000060000420004000000000000",
INIT_0F => X"0000024000240000102000000080000000000000000000240000800140000000",
INIT_10 => X"0080000000120CFC000000000000000001280013E010000000000900F8040000",
INIT_11 => X"2000000000000001480006D5801000000000000000091F0000800000004807C0",
INIT_12 => X"901A800080000000000000000820080006DD000000000000000002A00019DC00",
INIT_13 => X"0200800522C01252501086222082000010012024200000048019502000000C32",
INIT_14 => X"0080004501000200089400005200D0820008000000104C4800010600BC228404",
INIT_15 => X"0001040010000104001000010440080000822900000000801010500A13404111",
INIT_16 => X"32851951A0CA8080924C06403600086491900224002200400440104001040010",
INIT_17 => X"284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A128CA328CA",
INIT_18 => X"84A1284A1284A1284A1284A328CA328CA328CA328CA328CA328CA328CA328CA3",
INIT_19 => X"10000000000000000028CA328CA328CA328CA328CA328CA328CA1284A1284A12",
INIT_1A => X"69A69A250B61004055CD1439248209070CCCF48DE68A8900401038E2550A0010",
INIT_1B => X"341A0D068341A0D068A28A28A28A28A28A28A28A28A28A28A28A28A29A69A69A",
INIT_1C => X"56C1A0D269341A0D068349A4D068349A4D068341A0D269341A0D269341A0D068",
INIT_1D => X"0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE052",
INIT_1E => X"57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D00000000000000000000",
INIT_1F => X"D1575EF00557DF555D040000000043DF55087BC01EF007FD75FFFF84000AAFFD",
INIT_20 => X"7D5575455D557DFEF002AAAB55002E820AAAA843DFEF00517DEBA007BFDFEFFF",
INIT_21 => X"A28028AAAAAAABDF45F7803FFEF555568AAAF7802AA00FFFBD7555087BC00AAF",
INIT_22 => X"5087BD54BA550417400085155555082A95545552ABFE00087BC00AA082EBFE10",
INIT_23 => X"555D043DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00AA552E9554",
INIT_24 => X"BFFA2FBFFFFFAAD5400AAFF8402000A2FFFDF555D7BE8BFF5D51575EFA280175",
INIT_25 => X"000000000000000000000000000000000000000000557FF45002A975FF007BE8",
INIT_26 => X"D75D7FF84050BAEBDF78F45B68010482415B471C7E3DF451EFBEFBFAF4549000",
INIT_27 => X"17DE82007FFAFEFE3DB505EF1C5B7AF45490407000140038F450075C71FF087B",
INIT_28 => X"FFD55451C7FC70BAE3D155555415178FD7082EAAB550820870BAAA8438FFF005",
INIT_29 => X"07FC50BA002ABFE00AA8A2AABABEAEB8F45F78A3DFD741516DAAAE38E2DA28EB",
INIT_2A => X"FFFFC20BA5D2E905550071D54825D0A1543808515756D1C2497545552AB8E100",
INIT_2B => X"F5D55505FFBE801256D490E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92",
INIT_2C => X"451C24955EF0875EFBD7B6F1FFFC7BEDB45082EB8002000AAFFFDF6D417FEABE",
INIT_2D => X"5EFF7FBE8B5500000000000000000000000000000000000000000000000517DF",
INIT_2E => X"AB550055555FF007BD7555F784174AAA2FBEAB45F78402010007BD5545AAFFD5",
INIT_2F => X"174BAA68028BEF00517FE10007BE8BFFAAFFC01FF557FE8B550004174105D042",
INIT_30 => X"57FEAAAAAEBFEAAAAFFD5545557FD54BAAAD15754508556AB45002AA8B450800",
INIT_31 => X"04175555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7AAAAB45F7AEBFF45085",
INIT_32 => X"FD542000557FE8A00F3FFC00BA552E80145005557400552A954BA0051575EF55",
INIT_33 => X"A2FBFDFFF007FE8BFF5551401EFF784021FF002ABDFEFAAFBC00BA007BC0000F",
INIT_34 => X"000000000000517FF455D04155FF00557DF55FFD57DF55FFFBD5400A28400010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000004000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A14009801830084C182060000C10424840000000080000080200000000110204",
INIT_02 => X"0801080200100000046558040080000041000000002402400800000009008010",
INIT_03 => X"00020201040000D0842242024210810802006400088000003080054288C10000",
INIT_04 => X"0000400088020000003020002000001002A0E881108032100002000800203040",
INIT_05 => X"04092A081000411841480001000000201000012800400010001081C040402000",
INIT_06 => X"03600810100001220001E0001802002020240208000369001500100909000266",
INIT_07 => X"0000004000220440020000090C0810210A040004A0410000C0000810000C4901",
INIT_08 => X"0040480000802100100140004200808809000C002000000000010F8102041320",
INIT_09 => X"2008012000000000000200828888800808000410800840100220211850004442",
INIT_0A => X"040180240A80800442400004C0010000060210200008B2022304880800010000",
INIT_0B => X"0030000000010008008020020100008000400120800004004821202001A05A00",
INIT_0C => X"40510008101480000000A01004101480000000A0100000001300410402080080",
INIT_0D => X"0001A004101480000000A01004101480000000A0100540000040000000000000",
INIT_0E => X"00000000000040A8000900018040000000000000460800420004090000000000",
INIT_0F => X"0000034000082000102000000080028000000000000000240800800140000040",
INIT_10 => X"20900000001A00000002000000000020013000100010480000000D0000040440",
INIT_11 => X"2018000000000021500000800010440000000000400900008088000000680000",
INIT_12 => X"000000008200800000000000086010000080000100000000000082C000100000",
INIT_13 => X"000080000004924040008020000200101100004000000000C019500050000800",
INIT_14 => X"2B088A4541008240001000804000108280800001001051A12481041080801010",
INIT_15 => X"4480004800048004480044800044000240022100884000901210440003C14110",
INIT_16 => X"06E00000044200009849485D4020080000140004046240020044000480044800",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802000000400",
INIT_18 => X"0000000000000000000000020080200802008020080200802008020080200802",
INIT_19 => X"1000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"1451451AA654199951A24454514514F0CA940FE0D39712615FAD555204428290",
INIT_1B => X"CA6532994CA65329945145145145145145145145145145145145145145145145",
INIT_1C => X"670E572994CA6532994CAE572B95CA6532994CA6532B95CAE572994CA6532994",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE01C",
INIT_1E => X"03FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF0800000000000000000000",
INIT_1F => X"7FFDF45FFFBC2010AAD57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D0",
INIT_20 => X"0043DF55087BC01EF007FD75FFFF84000AAFF8002155AAFFE8B45AAD54000008",
INIT_21 => X"00557DF555D517FEBA082A801EFF7FBD5400FFD568B555D00155EF0804000000",
INIT_22 => X"AF7FBFDE00A2FBC0145005168A10AA843DFEF00517DEBA007BFDFEFFFD1575EF",
INIT_23 => X"EF5D7BC00AAF7D5575455D557DFEF002AAAB55002E820AAAA803FEBA082AAAAA",
INIT_24 => X"AAAF7802AA00FFFBD7555082E82155FFAEAAB55AAD568B455D00154BAFFFBD75",
INIT_25 => X"0000000000000000000000000000000000000000002ABDF45F7803FFEF555568",
INIT_26 => X"451EFBEFBFAF4549003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC700000",
INIT_27 => X"5EDB6DAADF470280075FFF45E3F1C7038A2DF78F45B68010482415B471C7E3DF",
INIT_28 => X"0A175C7000407000140038F450075C71FF087BD75D7FF84050BAEB8002155BEF",
INIT_29 => X"07FFAFEFE3DB505EF1C5B7AF45495B7DEAA0824851EFEBFBD2410EBD168B7D41",
INIT_2A => X"AA8038EAA0824A8AAAEBF5FAE28AAF1C2155005F68A10A28438FFF00517DE820",
INIT_2B => X"D4104104AAF7F1D75EF557FC70BAE3D155555415178FD7082EAAB550820870BA",
INIT_2C => X"45F78A3DFD741516DAAAE38E2DA28EBFFD55451C2087155EBA4A8B7DAADF68B7",
INIT_2D => X"FEFA2AEAAB55000000000000000000000000000000000000000000000002EB8F",
INIT_2E => X"2010007BD5545AAFFD55EFF7FBE8B5500043FE00F7D17FEBAA2D5574BAAAD17D",
INIT_2F => X"174AAA28002155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAB45F7840",
INIT_30 => X"BC2000AAD16ABFF002A975450004174105D042AB550055555FF007BD7555F784",
INIT_31 => X"8028BEF00517FE10007BE8BFFAAFFC01FF557FE8B55007FFDEAA0004175FFA2F",
INIT_32 => X"02AA8B450800174BAA68428AAA08042AABAAAD56AABAAAD140155087FEAA10A2",
INIT_33 => X"A2842ABEFAAFBE8BFF0004020AAFFD5555EF557FD54BAAAD15754508556AB450",
INIT_34 => X"0000000000002AAAB45F7AEBFF4508557FEAAAAAEBFEAAAAFFD5545550015555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000047FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B83008481800E0000C26426040000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"00080D4912E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"000048048002400048150000000002504230C899109032100020160880223000",
INIT_05 => X"040B2A229100410041088011100022201200012840440000B01088C0005C2400",
INIT_06 => X"03286A287E4003225021C5021880C02000A40249048363A5990010090908022A",
INIT_07 => X"8320694044222987020C80152D8910210A0400252B74200045C86810000C5B05",
INIT_08 => X"00404126509804400501400242C0B0B83B0134702000000000191FA162841324",
INIT_09 => X"2008013002000220001240820F8B2A08000040409018401001200159D80D64AA",
INIT_0A => X"91019B02080885200042E098C00101B0070310200008B60A23A51B2802067327",
INIT_0B => X"003000080802500C088325828102408120409120940680100504022148504440",
INIT_0C => X"1501D5761B011986695014A96E1A8119865A5018C5A0A00012004104020808B0",
INIT_0D => X"A2600AAE1A811986695014A96E1B0119865A5018C5AF0062C38A4DB680A0D824",
INIT_0E => X"1DB528802CAB184E8F4101621B1BAC845542056A289A1BB2078A922DA2A8B180",
INIT_0F => X"7A3D94392000224ACDE215883078681B5C05AA429189B60AC43CEC7F0272C384",
INIT_10 => X"134CD551BCA1C90006C0C2958502861120C003104289A668B8CAB27010633831",
INIT_11 => X"82806CA64090B89E015AAA880E48382EB8804B020A06020C67061BC785938085",
INIT_12 => X"470126C6284B2D20410AB4503089C00A8280819A5539D503336D61056ABA0062",
INIT_13 => X"000080060040142020015001004A00080042004000E8089C9003066E03513E41",
INIT_14 => X"010CBA45367082014000908020349320008000A1000C09A9348498B000000000",
INIT_15 => X"C32A0832A0C32A0C32A0832A0C19504195040040000000801010028001400010",
INIT_16 => X"2468118104400000904C0C0964200841010954000444D280140050C32A0832A0",
INIT_17 => X"4090240902409024090240902409024090240902409024090240902409024090",
INIT_18 => X"0100401004010040100401024090240902409024090240902409024090240902",
INIT_19 => X"0000000000000000004010040100401004010040100401004010040100401004",
INIT_1A => X"410410502A441495418984700000005088804180C0B10A04D0A7104201400284",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000010410410",
INIT_1C => X"7800000000000000201000000000000000000008040000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE060",
INIT_1E => X"4155EFAA842ABEFA280155EFFFFBC01EF0855400005500000000000000000000",
INIT_1F => X"FBFFF4508514000000003FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF080",
INIT_20 => X"280154BA5555401EFFFD5421EFA2FFFFF555D51575FFA2FFD75FF550015400FF",
INIT_21 => X"FFFBC2010AAD568AAAAAD142145FF80155EF0051555FF0804155FFF7D57DF45A",
INIT_22 => X"008001540008514215555003DFFFA28002155AAFFE8B45AAD540000087FFDF45",
INIT_23 => X"0000040000000043DF55087BC01EF007FD75FFFF84000AAFF802ABFFA2AABFE1",
INIT_24 => X"400FFD568B555D00155EF085168B45085142010FFAE800AA5D7BFDF45F7FFEAA",
INIT_25 => X"000000000000000000000000000000000000000000517FEBA082A801EFF7FBD5",
INIT_26 => X"7DF7DA2AEB8FC70000175EFB6802DBC7BE8A155EFE3FBC71FF145B4203855000",
INIT_27 => X"5D05EF550E15400E3F1FFF7D085B420381C003DE10BEF5EDAAAAAD547038EBD5",
INIT_28 => X"04105C7F7DF78F45B68010482415B471C7E3DF451EFBEFBFAF45495F575FFBEF",
INIT_29 => X"ADF470280075FFF45E3F1C7038A2DB68ABAB6D145145FF84155D7085B555C714",
INIT_2A => X"EB8428BEFBEA4BDE28140A1543800514515549003FFC7BE8002155BEF5EDB6DA",
INIT_2B => X"2417FFFF7DE3F1EFA10140407000140038F450075C71FF087BD75D7FF84050BA",
INIT_2C => X"AA0824851EFEBFBD2410EBD168B7D410A175C7005B6DB55145140000FFAE8508",
INIT_2D => X"5EF557BC20AA5D0000000000000000000000000000000000000000000005B7DE",
INIT_2E => X"FEBAA2D5574BAAAD17DFEFA2AEAAB550004175FFF7803DF45FFAE955EFAAFBD5",
INIT_2F => X"E8B55007FD75FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D043FE00F7D17",
INIT_30 => X"015555007FD5545550400145FFFBEAB45F78402010007BD5545AAFFD55EFF7FB",
INIT_31 => X"8002155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAAAAFFD555545FF8",
INIT_32 => X"07BD7555F784174AAA2842ABEFFF803DEAA5D2E974AA00515754500003FF55FF",
INIT_33 => X"555540000FFAE97410007BFFFFFA2D57FE105D04174105D042AB550055555FF0",
INIT_34 => X"0000000000007FFDEAA0004175FFA2FBC2000AAD16ABFF002A97545007FFFF45",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000004000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C048000C048400380000007024040000000080000088200002802153231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"421A0A0012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"02004000890200001837800001998C31C090609C104000102002140900003548",
INIT_05 => X"0402002BC200009841090001200006200800000020480010A4100100001C2000",
INIT_06 => X"033432287FC003230001D0001806C0060CB0622000037085C800100C0C200008",
INIT_07 => X"135038CE64B663DFA314C803292140890C0601F472D1640051F80C10020C493F",
INIT_08 => X"00000167C081000011814004C20481A92940EA7A3020480000071F846890162E",
INIT_09 => X"D40C01240008000080024082488BAF08000020000208401004300421800F04F8",
INIT_0A => X"F9F80FA0200E0BF40063FF9DC0010000180018200408B27E234913E900067F04",
INIT_0B => X"001100002002801000A04200000000000000000000029D204B7C0382FD0100F3",
INIT_0C => X"9628F97E0B348EDAC3900F6EFA0B158EDA93900F6EE230381208008001007A80",
INIT_0D => X"EAE64BCA0B158EDAC3900F6EFA0B348EDA93900F6EE8421392C96B1237E0D8BD",
INIT_0E => X"4CAEAD412EDD2B47CFF812A383430C669E622DBC31D73F6006A5891533EF9500",
INIT_0F => X"2E19B8BA30E022DAD8C100CA39E8CEBE66C2B083798D341B10DE7E14400392C7",
INIT_10 => X"32966471A9C5DD00B12728D5360234D62A49FAB442994B3238D4E2FB10463665",
INIT_11 => X"F0FABAC800DA550C29F36A8A2554E48A6430469392526208C6CC95C33717D885",
INIT_12 => X"2B416A51B60585A5C28895962502E9F36A828C4999AF580395542D27CDBA0020",
INIT_13 => X"0000800000001E404011F066000A000EE040000000873FB80B8A00EF03F56CC1",
INIT_14 => X"2284304D667C06CC6816B300403C13E2000000460010400000010CE080801010",
INIT_15 => X"872F0872F0C72F0872F0872F0C597863978421000800209010104ACA03414110",
INIT_16 => X"01000000104280009048004000000800001D5E05182493C5BC5AF0872F0C72F0",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0802008020080200802008000000000000000000000000000000000000000000",
INIT_19 => X"1000000000000000000080200802008020080200802008020080200802008020",
INIT_1A => X"492492240F010000146E502D4514510246088881360A95118B120CB054420210",
INIT_1B => X"6432190C86432190C82082082082082082082082082082082082082092492492",
INIT_1C => X"7FEB2592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2590C8",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"5421FF00042ABEFFF8400010082EAABFF55002ABEF0800000000000000000000",
INIT_1F => X"002ABEFFFFBD54000004155EFAA842ABEFA280155EFFFFBC01EF085540000555",
INIT_20 => X"AFBE8AAAA2D540000F7D57DF55A2AABFFEF08556AA10000028AAAFFD15541000",
INIT_21 => X"085140000005168AAA087BFFFFF5D04001FF00041554555557FE005D003FE10A",
INIT_22 => X"F0851555FF082AA8B55F7AEA8BEF5551575FFA2FFD75FF550015400FFFBFFF45",
INIT_23 => X"10AAD57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D0000145082E955F",
INIT_24 => X"5EF0051555FF0804155FFF7842AA100000020BAAA801541055042ABEFFFFBD54",
INIT_25 => X"0000000000000000000000000000000000000000005568AAAAAD142145FF8015",
INIT_26 => X"C71FF145B42038555F401D71C0A2DBC7EB80000280824ADBD7490E28BEF08000",
INIT_27 => X"A2DA82FFDB5243800002FBD7EBFBD24101C00175EFB6802DBC7BE8A155EFE3FB",
INIT_28 => X"5B7AE1041003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7005F6AA381C0",
INIT_29 => X"50E15400E3F1FFF7D085B420381C5B6AA82147FF8FEF410E001FF000E1755555",
INIT_2A => X"49000017D142E905EF1451525C7082AADB45F7AEA8BEF555F575FFBEF5D05EF5",
INIT_2B => X"041002FBEFEBFBD2410AADF78F45B68010482415B471C7E3DF451EFBEFBFAF45",
INIT_2C => X"BAB6D145145FF84155D7085B555C71404105C7F7842FA381C0A00082AA8A1041",
INIT_2D => X"F55002AA8BEF000000000000000000000000000000000000000000000005B68A",
INIT_2E => X"DF45FFAE955EFAAFBD55EF557BC20AA5D7BC01555D2EBFF55A284000AA08003F",
INIT_2F => X"AAB55007BE8AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D04175FFF7803",
INIT_30 => X"E821FF082A97555557FE8A0000043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AE",
INIT_31 => X"7FD75FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D7BE8A005D7FEABFF002",
INIT_32 => X"AFFD55EFF7FBE8B550004001FF5D2A801EF5D5142145082EBFF55F7AAAABEF5D",
INIT_33 => X"552A82010A2AA8000008043FFFFA2FBC2010A2FBEAB45F78402010007BD5545A",
INIT_34 => X"0000000000007BEAAAAFFD555545FF8015555007FD5545550400145FF843DEAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400986B830E84D182260000C1042684001000008220008A20019080A510200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00020201926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"00104884880A4400403003005800027102A0E8C110D83210642EA809C0203040",
INIT_05 => X"04092A08138041184109C001380000201A008128044E00754010C9C192D82400",
INIT_06 => X"032C7E201800012372A1D72A180000204024024954A3670819001009092C0222",
INIT_07 => X"0164004000220B40020C80052C0A12292A040005715540015E006810001C4B01",
INIT_08 => X"0040549032881001140140024200808839005C002010800000155F8122851320",
INIT_09 => X"6008012C80481284881280825A988008000040808629441005B3071859006442",
INIT_0A => X"0001B0200810940400720005C0030192072310200028B6022346080802E001A5",
INIT_0B => X"003000206822F20CA8826AC2A14250A128509528954404144C20042501004000",
INIT_0C => X"03D404A41AA5B7344C10B383081BA4B7341C10B3831034081200000000000430",
INIT_0D => X"5A2B2C381BA4B7344C10B383081AA5B7341C10B383110218CB0E54C2EA404A4F",
INIT_0E => X"3548B3A008E730A01AB113A5524E6ACA678001CE3E20A5B284ED1132909C7288",
INIT_0F => X"0A3C066430202021252991C22C99731014AC3CC0C0B8182597A801610218CB0C",
INIT_10 => X"A5C8825194332B018A444AEA2701288A15A151EC5952E44128CA194517354C18",
INIT_11 => X"635232D50048A411C158BB0A7910142C771804C8A0ADA2E6A983014780CA28B2",
INIT_12 => X"6E4023F8BE8E3E1E0109472C3EB50158BB02D09852745F80112C428562EE0353",
INIT_13 => X"00008002414032646000826080C20001104240480068001C9B9150A000029704",
INIT_14 => X"1118BA4510008241C80290882400908000A000A1000809A93485D61000000000",
INIT_15 => X"40000000000000040000000000000020000000040000008010122A8201410058",
INIT_16 => X"246A10A1044101A89A4D0C096420184321040002844840000000004000000000",
INIT_17 => X"5094250942509425094250942509425094250942509425094250942509425094",
INIT_18 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_19 => X"0000000000000000005094250942509425094250942509425094250942509425",
INIT_1A => X"75D75D7FEDFDFDFDFBEEF9DD555555F7EEFF3F7DF7FF3E7E1FBF7DF7E24502A8",
INIT_1B => X"FAFD7EBF5FAFD7EBF5D75D75D75D75D75D75D75D75D75D75D75D75D75D75D75D",
INIT_1C => X"7FEFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F780000000000000000000",
INIT_1F => X"AA97400AAD540155A2D5421FF00042ABEFFF8400010082EAABFF55002ABEF085",
INIT_20 => X"A842ABEFA280155EFFFFBC01EF08554000055043DEBAF7843FFFFF7AABDF55A2",
INIT_21 => X"FFFBD5400005568A1055043DEBAAAFFE8B45557FD7410552EAAABAAA84155EFA",
INIT_22 => X"AA2FFE8ABAAA8428A00087BD7555FFD56AA10000028AAAFFD15541000002ABEF",
INIT_23 => X"55A2803FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF085557545FFD17DEB",
INIT_24 => X"1FF00041554555557FE005D0000155557BEAABA5D2ABDF450851420AA5D7FD55",
INIT_25 => X"0000000000000000000000000000000000000000005168AAA087BFFFFF5D0400",
INIT_26 => X"ADBD7490E28BEF08516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EB800",
INIT_27 => X"03FFD7EBA4BDF45AAAA90410BEDF45155A2DF401D71C0A2DBC7EB80000280824",
INIT_28 => X"2AAFA82B680175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550E38E92EB8",
INIT_29 => X"FDB5243800002FBD7EBFBD24101C556FA38490A3FE92BEFFEAB45417FD24385D",
INIT_2A => X"00515056DE3D17FE92BEF1EFA92AA8428A10007FD557DFFDF6AA381C0A2DA82F",
INIT_2B => X"5085B400925D7FD557DA2803DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7",
INIT_2C => X"82147FF8FEF410E001FF000E17555555B7AE10410E00155497FEFABA4120B8F5",
INIT_2D => X"ABAA2FBD7545AA8000000000000000000000000000000000000000000005B6AA",
INIT_2E => X"FF55A284000AA08003FF55002AA8BEF00517FE00082EBDF45AA8428A10085568",
INIT_2F => X"C20AA5D2EA8A00A2803DF45AA843DF55AAAE82000F7FBD5545AAFBC01555D2EB",
INIT_30 => X"FE8B55087FC00BA552ABFE10F784175FFF7803DF45FFAE955EFAAFBD55EF557B",
INIT_31 => X"FBE8AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D517FEAA082EBFE10F7F",
INIT_32 => X"AD17DFEFA2AEAAB550051401FFA2D57FE10F7D57DE00AA842AA00007FD75FFF7",
INIT_33 => X"007BFDEAA08042AB45087FC0010557FD55FFAA843FE00F7D17FEBAA2D5574BAA",
INIT_34 => X"0000000000007BE8A005D7FEABFF002E821FF082A97555557FE8A00002E82155",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000067FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"0002074F200904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000480488024000403000000000001002A0E881108032100002000800203040",
INIT_05 => X"04092A081000411841080001000000201000012800400010001081C000402000",
INIT_06 => X"033D7880500001221021C1021800002000240249048361001100100909000222",
INIT_07 => X"9020304000220050020480152D0A142D0A8400043B45400040006810000C5901",
INIT_08 => X"0040400010880000100140024280808829029C002000000000053FA142051324",
INIT_09 => X"6008012000000000000200820888800800004000800840100020011858006442",
INIT_0A => X"000110200800840400400005C0010190070310200008B202236D080802000001",
INIT_0B => X"003000000000100C088020028102408120409120940404104C20002101004000",
INIT_0C => X"2050805210040000B0E0A0000210040000E0E0A0000190081200000000000000",
INIT_0D => X"0111300210008000B0E0A0000210008000E0E0A0000B02740421A0E5D1A02400",
INIT_0E => X"C0715C40110080A4006110510C14D18178E01200860008920106460D4501CB00",
INIT_0F => X"500002411420220080220C0093C38923240ABBC00905C33C6000400F02740412",
INIT_10 => X"9682398000120800658992F3C700C3018120000041DB011CC000090012565306",
INIT_11 => X"B7A0B1E240240A8340000200067EAA8CB65809240C09024A4AE0CA0000480083",
INIT_12 => X"00845C7DB0D0200900422ACA4B28000002002B46867DBC002A830280000800F7",
INIT_13 => X"000080020040126060008020000200000042004005800004801150A003412440",
INIT_14 => X"01088A4500008240000000802000908000800001000009A92481041000000000",
INIT_15 => X"0000000000400000000000000400000000000000000000801010000001410010",
INIT_16 => X"246810810440000090480C096420084101040000044040000000004000040000",
INIT_17 => X"4090240902409024090240902409024090240902409024090240902409024090",
INIT_18 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_19 => X"0000000000000000004090240902409024090240902409024090240902409024",
INIT_1A => X"3CF3CF3FE77DDDDD55E6D5FCF3CF3DF7CE5C8FF0F7BE9D75CF9F7DF650400280",
INIT_1B => X"FE7F3F9FCFE7F3F9FCF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"8007F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE07F",
INIT_1E => X"17DF45AAD157400007BEAAAAAAAE955555D5568A105D00000000000000000000",
INIT_1F => X"AA800AAF784020AAF7D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7D",
INIT_20 => X"0042ABEFFF8400010082EAABFF55002ABEF085155400FFD1420100055574AAA2",
INIT_21 => X"AAD540155A28028B550051574005D7FFFE105D7BD7545A284020BA0055421FF0",
INIT_22 => X"00851421FF5D7FFDEBA085168B45FF843DEBAF7843FFFFF7AABDF55A2AA97400",
INIT_23 => X"FF5504155EFAA842ABEFA280155EFFFFBC01EF08554000055002AB455D514201",
INIT_24 => X"B45557FD7410552EAAABAAA8017400AAD140000002EBFFEFA2AAA8BEFF780021",
INIT_25 => X"0000000000000000000000000000000000000000005568A1055043DEBAAAFFE8",
INIT_26 => X"F8E38E3DF45155EBD17FF6DAADB504001C71EDA82AAA0955455D556DA0049000",
INIT_27 => X"B420101C55554AAAAA480082FF84000BAEBD16DA82410A3FFD7AAA4B8E824971",
INIT_28 => X"8405092085F401D71C0A2DBC7EB80000280824ADBD7490E28BEF085157428FFD",
INIT_29 => X"BA4BDF45AAAA90410BEDF45155A28E2AB7D0051504005D71F8E004975D556DB6",
INIT_2A => X"550028B6D5D51420101C5B401EF417BFAEAA08516AB45E38E38E92EB803FFD7E",
INIT_2B => X"7A2AEAFBC7EB80071FF5500175EFB6802DBC7BE8A155EFE3FBC71FF145B42038",
INIT_2C => X"38490A3FE92BEFFEAB45417FD24385D2AAFA82B68015400AADB40000082EBFFC",
INIT_2D => X"54555557FE1000000000000000000000000000000000000000000000000556FA",
INIT_2E => X"DF45AA8428A10085568ABAA2FBD7545AAD17DFFFAAFFC200055557DE00A28015",
INIT_2F => X"A8BEF0051554AAFFFFC00105D55554BAA28400000F784020BAAAD17FE00082EB",
INIT_30 => X"568A000051575FFF78415410087BC01555D2EBFF55A284000AA08003FF55002A",
INIT_31 => X"AEA8A00A2803DF45AA843DF55AAAE82000F7FBD5545AAAEAABFF0051400105D5",
INIT_32 => X"AFBD55EF557BC20AA5D042ABFF555142000557FC01EF007FEAABA00556AB55A2",
INIT_33 => X"A2FBC0010082EBDF55A2AABDF45A284175FF5D04175FFF7803DF45FFAE955EFA",
INIT_34 => X"000000000000517FEAA082EBFE10F7FFE8B55087FC00BA552ABFE10F78415400",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000100000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"000440009282000001100000000000100220C8811080321000000228002A3000",
INIT_05 => X"04092A0010004300418800510000A6201000012A64400000145080C000422000",
INIT_06 => X"032B1800100001220001C00018821020402402080003772019001009090002AA",
INIT_07 => X"0000004000220000021840010C8912250A0400042044400040006810000C4901",
INIT_08 => X"0040400022810000058140024280A0A8190004002030C00000016F8122041320",
INIT_09 => X"E0080120000000000002C0820888008800000000800840100020011850004402",
INIT_0A => X"00013000080094000062000180010180060210200008B2022304080800000003",
INIT_0B => X"0030000000000008008020020000000000000100800000000000002500004000",
INIT_0C => X"0000000010108000000000000010108000000000000230001200000000000420",
INIT_0D => X"0000000010140000000000000010140000000000000100000040000000000000",
INIT_0E => X"0000000000000000000100008040000000000000000000020000090000000000",
INIT_0F => X"0000000030002000406000000000068409014000000000000000000100000040",
INIT_10 => X"2010000000000800000201000800000000000000400048000000000010000440",
INIT_11 => X"00184400A0000000000002000000441108800000000002008008000000000080",
INIT_12 => X"0000000242038B82800000000000000002000001000000000000000000080000",
INIT_13 => X"000080000000100000000005C04A000000400000000000000001062000000400",
INIT_14 => X"01088A4500008200000000800000100000800001000001A12480001000000000",
INIT_15 => X"4000040000000000000000000400002000020000000000801010000041400010",
INIT_16 => X"0460000004400000904808094020080000000000044040000000004000040000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000400280",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FC00000804154AA5D00001EFF78428AAA007BC2145F780000000000000000000",
INIT_1F => X"55400AA007FC2000F7D17DF45AAD157400007BEAAAAAAAE955555D5568A105D7",
INIT_20 => X"D043FFFFAAAABDEAA557BFDE00FFD140155F7FBD74AAAAD17DF45F7D1421EF00",
INIT_21 => X"F784020AAF7FFFDF45FF84000BA552ABDFEF08517DF55A2FBEAB555D556AAAA5",
INIT_22 => X"5AAFFEAB45F7843FF45082A801FF005155400FFD1420100055574AAA2AA800AA",
INIT_23 => X"AAA2D5421FF00042ABEFFF8400010082EAABFF55002ABEF087BE8ABA555168B5",
INIT_24 => X"E105D7BD7545A284020BA007FFFE10A284000AA0055401550055574005D2E800",
INIT_25 => X"0000000000000000000000000000000000000000000028B550051574005D7FFF",
INIT_26 => X"955455D556DA004971C7038140012482550E021C7EB8028A821C7BC516DFF800",
INIT_27 => X"17FF45E3DF471C70851400BA0071C5028FFD17FF6DAADB504001C71EDA82AAA0",
INIT_28 => X"FBE8B555D516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBF1D5492BED",
INIT_29 => X"C55554AAAAA480082FF84000BAEBF1FFF7DEB8000092552ABFFEF08517DF6DB6",
INIT_2A => X"087FEFA8241516DB55A2FFEAB6DEB843DF551C20801C71C5157428FFDB420101",
INIT_2B => X"5085550428412A85082BEDF401D71C0A2DBC7EB80000280824ADBD7490E28BEF",
INIT_2C => X"7D0051504005D71F8E004975D556DB68405092087FF8E00BE8A02082005F4714",
INIT_2D => X"A00557BD75EFF78000000000000000000000000000000000000000000000E2AB",
INIT_2E => X"200055557DE00A2801554555557FE100055554BA5504000105D2A80145AA842A",
INIT_2F => X"D7545AAD557410F7D57DF55AAFBD55450055420BA0055574BAF7D17DFFFAAFFC",
INIT_30 => X"ABDFFF08517FFFFF7FBEAB455D517FE00082EBDF45AA8428A10085568ABAA2FB",
INIT_31 => X"51554AAFFFFC00105D55554BAA28400000F784020BAAAD57FFEFA28402010552",
INIT_32 => X"8003FF55002AA8BEF007FFDE1000557DF45AAFBE8BEFA2803FF4555040015555",
INIT_33 => X"F7AE80000087BD55450855400BA002A95400F7FBC01555D2EBFF55A284000AA0",
INIT_34 => X"0000000000002EAABFF0051400105D5568A000051575FFF78415410087FEAA10",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000006000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"0202115002BB10080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"2FE962000017102918900948514522CE09200C0D590569398ADBF8CC1E50E480",
INIT_05 => X"5E6023002834854AE41C1E8782F508F2A15B71D412E0AFD9C2990DA56FF0B55A",
INIT_06 => X"82A803B9B9E55402000340003200220A86012D0000000480D02A7960540180A0",
INIT_07 => X"01380C40D890101DBD400901442800817C2901F400868554DE240000A80090CE",
INIT_08 => X"18A9050122004000005665510320C9C90510025A8A00000A0A048F550A440E00",
INIT_09 => X"2A8A562060410280081116C8204D016CB2CB2900080082795804112890000001",
INIT_0A => X"4052E400008176802200020025699200140001A15000017F0051D0F837324E00",
INIT_0B => X"5514554485D000000124002400000000000001004010A8812831605DA0000A05",
INIT_0C => X"708E2CB5320018CAC99BA0A3B9320018CAAAADA0C343F1AC1B01040A00202489",
INIT_0D => X"E7A3EE59320018CAC99BA0ACB9320018CAAAADA0CC421CA003B694B68018FAAA",
INIT_0E => X"24352AB2449A3FF2FA04E5E09B128834ADB1443A1891E4A928C29020E6A8524C",
INIT_0F => X"714C902375B801324301AB0067622E5E5404B2A5A40B1E6644AF0F021EA003AC",
INIT_10 => X"1216F50A8C241815FEB6A9158863F638FB60ED838E890B703C6260D8E3A21275",
INIT_11 => X"555E4C15F11133D171727A2550EE2F1BA0064F70DBDB1C74424E91E1C194C71D",
INIT_12 => X"ACCC59432A2B2D001F803471A9A960E57245FDF9D364DBD9435A6D45C9E81BED",
INIT_13 => X"0012CAC00006B0800000038814B72AB01508150013F162119014204373517700",
INIT_14 => X"002912300208092B940192D1000000000000A8A5AA80018120E0006600000000",
INIT_15 => X"1100011000110001100011000108000880008000520228080108039501200848",
INIT_16 => X"012000081500008A422150884081AC9000010003561180063DB4F61100011000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"28A28A3D2DE5F87963445469E79E7853D44C690DA64C1C69818768A360400000",
INIT_1B => X"F4FA3D3E8F4FA3D3E9A29A29A29A29A29A29A29A29A29A29A29A29A28A28A28A",
INIT_1C => X"000FA7D3E9F4FA7D1E8F47A3D1E8F47A3D1E8F4FA7D3E9F4FA7D3E9F4FA7D3E8",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"43FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE005500000000000000000000",
INIT_1F => X"80020005D2A95410FFFFC00000804154AA5D00001EFF78428AAA007BC2145F78",
INIT_20 => X"AD157400007BEAAAAAAAE955555D5568A105D2E974BAF7FBEAB45FFFFC00BAF7",
INIT_21 => X"007FC2000F78000010552E800AA002E821FFA2AAAAA00000417555FFD17DF45A",
INIT_22 => X"A08043FEBA5D55575FFF7AABFE00557BD74AAAAD17DF45F7D1421EF0055400AA",
INIT_23 => X"10FFD56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7AABDF55F7AE820A",
INIT_24 => X"FEF08517DF55A2FBEAB555D04154BAA2FBE8B55FFFFD55FF557FC2000FF80154",
INIT_25 => X"0000000000000000000000000000000000000000007FFDF45FF84000BA552ABD",
INIT_26 => X"28A821C7BC516DFF8438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE1049000",
INIT_27 => X"BE8B55FFF1C70BAF78A000005D2097438FFF1C7038140012482550E021C7EB80",
INIT_28 => X"0E1757DEBD17FF6DAADB504001C71EDA82AAA0955455D556DA00492490492F7F",
INIT_29 => X"3DF471C70851400BA0071C5028FF84020285D2085092002A801FFB6AAA8A1008",
INIT_2A => X"EBA4BAF6DE3AA8709208043FEBA555B555FFE3AABFE005D71D5492BED17FF45E",
INIT_2B => X"7557BC0028E38412428EBD16DA82410A3FFD7AAA4B8E824971F8E38E3DF45155",
INIT_2C => X"7DEB8000092552ABFFEF08517DF6DB6FBE8B555D04124BAB6FBE8B45E3FBD55D",
INIT_2D => X"55555003DE000000000000000000000000000000000000000000000000071FFF",
INIT_2E => X"00105D2A80145AA842AA00557BD75EFF78428B55AAD168B55F7FFFDFEFFFAA95",
INIT_2F => X"7FE10000000010F7FBEAB45FFD1554AAFFAE820105500154AAF7D5554BA55040",
INIT_30 => X"E801EFF7AEA8A10002E955FFA2D17DFFFAAFFC200055557DE00A280155455555",
INIT_31 => X"5557410F7D57DF55AAFBD55450055420BA0055574BAF784000BA5D0017410082",
INIT_32 => X"85568ABAA2FBD7545AA802ABEFA2AA9541000003DEBA557BD75EFA2AEBDE105D",
INIT_33 => X"FFFBEAB45AAFFD55555D7FC20AAA280000AAAAD17FE00082EBDF45AA8428A100",
INIT_34 => X"000000000000557FFEFA28402010552ABDFFF08517FFFFF7FBEAB455D04020AA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000002000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"5295B6957FCBE0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"6DE90201BF90102103AF158E805428249851BFB2C106592088DBF8400A5055C2",
INIT_05 => X"3824BD7F80148D9E07100A8201ED01C1A19B68F40A807ED9C18114956FF081DB",
INIT_06 => X"ED08CA6A8F033DD800000000050716BE9F57F8AC000807DFD999E0E5E1818B1B",
INIT_07 => X"00150886481240FE05A109228E2C0891D772A6F40045B8CF30E085DD2ED57D4E",
INIT_08 => X"72637FDF23800005981C0338190549C904182B6113870022000488C08B46268A",
INIT_09 => X"3E7437823DF78CDB6CA60E0E28EFFE2061872F80C1684A80C8604085F0074D3B",
INIT_0A => X"F5B4FFBD2FAD7FE653C36A1FF33E0E001E000B3A5DAADAFDDA5DA79350CFB801",
INIT_0B => X"CFE833C5C3D00018006C681700000000000000020012E9E10A31EB5FF9296A67",
INIT_0C => X"0D5ECE542A6FEEB2533EA160782A6FEEB2333EA16031F2BD47BDA2CA5D8164FC",
INIT_0D => X"282400F82A6FEEB2533EA160782A6FEEB2333EA160391BEFF2C32FB695F91911",
INIT_0E => X"573FAD5A86840354D1706FFFA3EF6E24B6D18C0D06638A207CFDE1F7DDAD76D5",
INIT_0F => X"FE4ACA4D77FAAB77CE3AF3EE78F58DB737E6E43E59AFE4A59B57679D19EFF2C7",
INIT_10 => X"ADB55572CA52606DFED6CA55334C04C04FF7D7A0ABD6DAAAB96529382B74E4E1",
INIT_11 => X"F9956EAA1A184045D5D7A870D2F5A5D7522D1281017F056E9C9C3FC95949C157",
INIT_12 => X"1F432EA58949D5B5C85F97871876F7D7E859FDEB974F486905001FDF5FA0D719",
INIT_13 => X"DEF20670021EE341036BF368128419FB5560158015177F916A039EF41FDB34A9",
INIT_14 => X"00633F1D0A7CC9AE7A08BFF0001D35682AC0CE8FCCC200A59BDD2FFE3F3EC7C7",
INIT_15 => X"FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A7800617112E46F05D02DD814102F8",
INIT_16 => X"05F08000179C16DECF67F08BC02F9086000D9E8A3F06ABD73DBCF4FBCF4FBCF4",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"34D34D48C4986868DC800181D75D7445F009EDCC4052E92E0204114F981800C0",
INIT_1B => X"1A8D468341A8D46834D35D74D34D35D74D35D74D34D35D74D35D74D34D34D34D",
INIT_1C => X"0008D46A351A8D46A351A8D46A351A8D46A351A0D068341A0D068341A0D06834",
INIT_1D => X"0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"43FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF5500000000000000000000",
INIT_1F => X"8028A00F7843FEBA55043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE00550",
INIT_20 => X"804154AA5D00001EFF78428AAA007BC2145F7D568B45000002010552EBDF45A2",
INIT_21 => X"5D2A95410FFAE800105D2A95410002A95410AAAEBFF55AAFFC00BAF7FFC00000",
INIT_22 => X"FFFD57DE00F7AE800AAAAAABDFEF5D2E974BAF7FBEAB45FFFFC00BAF78002000",
INIT_23 => X"AA5D517DF45AAD157400007BEAAAAAAAE955555D5568A105D7FFFFEFA2D568BF",
INIT_24 => X"1FFA2AAAAA00000417555FF8028B55082A974105D003FF55F7802AAAAAAD168A",
INIT_25 => X"0000000000000000000000000000000000000000000000010552E800AA002E82",
INIT_26 => X"955C71C043FE10490A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD749000",
INIT_27 => X"E050384124BFF7DB68A28A38F7803DE82490438FC7E3F1EAB55B6DF6DBFFF7AA",
INIT_28 => X"F5C70BAFFF1C7038140012482550E021C7EB8028A821C7BC516DFFDF68B551C0",
INIT_29 => X"FF1C70BAF78A000005D2097438FFAA85000492495428082E95400AAA0BDF7DB6",
INIT_2A => X"497FFAFFFB6D56FBFFEBDB78E38F7AA800BAB6AEBDFD75D2490492F7FBE8B55F",
INIT_2B => X"DEB8028AAAB6D16FA8249517FF6DAADB504001C71EDA82AAA0955455D556DA00",
INIT_2C => X"285D2085092002A801FFB6AAA8A10080E1757DEB8A2DB5514249243841003FF6",
INIT_2D => X"0BAF7FFFDF550000000000000000000000000000000000000000000000004020",
INIT_2E => X"8B55F7FFFDFEFFFAA9555555003DE00002ABFFEFF7FBFDFFFAAD168B55AA8000",
INIT_2F => X"D75EFF7FBEAB45552E954BA08003DFFFFFAAA8AAAF7843FE10000428B55AAD16",
INIT_30 => X"E95410AA843FFFFF7D5554BAF7D5554BA5504000105D2A80145AA842AA00557B",
INIT_31 => X"0000010F7FBEAB45FFD1554AAFFAE820105500154AAF7AE974000800154AA002",
INIT_32 => X"2801554555557FE10007FEABEFFFD57FFEFAAFFE8ABAFFAA820BAF7AEBFF5555",
INIT_33 => X"5500020AA08003DFFFA28028AAAF7D17DE0000517DFFFAAFFC200055557DE00A",
INIT_34 => X"00000000000004000BA5D0017410082E801EFF7AEA8A10002E955FFA2AABFF45",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000067FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"080BA868803F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"42016B0C401F58495C900A4859552A611D9A640F5903B2388004004C08A06008",
INIT_05 => X"16226B107811422A641C08038040007060E0032801E0202000991B708280B501",
INIT_06 => X"120886B3B8E0FC86142B4142B0000000011114D3058240240907F82000000000",
INIT_07 => X"006880802102401015610A02C4005000EA019D002482043FCF1C8090C02800C0",
INIT_08 => X"11018020D40A5004003260F9810541494D403D9B98810A0002C601000054B94A",
INIT_09 => X"022E0C6070000504102805C820C8016C30C250080C0182183804012A0A102200",
INIT_0A => X"084001E000108010230495A800FD865421432121804021C20452880C2D100000",
INIT_0B => X"3F140FC2060014250B9080008306C18360C1B0609C05013065CC042004040808",
INIT_0C => X"DF7C728582081483ACC15F9C3982081483CCC15F9CBA45505640000A40201900",
INIT_0D => X"DFEBFBF982081483ACC15F9F3982081483CCC15F9FB1962FCB69E08AAAEAEBCD",
INIT_0E => X"CAA02FE3F8E7F5E3AC3620805298B15A3FEBF1CFFF7670ACC3811A28AB57523C",
INIT_0F => X"01BD67DC4041D4CF03138DD865103EFEEAC9002BF05800D875E63CC9962FCB52",
INIT_10 => X"0016EA8DB7BFE25208E8F46A228BF8A757F1B72A8A800B7546DB9F1CA320037F",
INIT_11 => X"81A8A29509EAAE7FD3B749471C48F8A45981CCFAFDBF9464006FD037AEFAE515",
INIT_12 => X"EFF5778802A3AF8E8FB0440CE78773B709641256EC844B8AF92FD7CEDC24A9E1",
INIT_13 => X"0003C1C284601C2864000080113307E4800297D086E00036D2440E0880AAD62B",
INIT_14 => X"C44C92A88DCC2211E44174112840880000060D7030C30B885200D27400400808",
INIT_15 => X"0030800308003080030800308001840018400400602A01880980037109700C04",
INIT_16 => X"6808348340000020301805002D008CD943626111C0D95C20C2030A0030800308",
INIT_17 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B0",
INIT_18 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_19 => X"00000000000000000041B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_1A => X"1451451223059150A2EFB05C104104B3CEB80EE173C2300FCA8B7DF160000000",
INIT_1B => X"4AA552A954A25128955545145145155555545145145155555545145145145145",
INIT_1C => X"00025128944A25128944A25128944A25128944A25128944A25128944A2512894",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"43FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA0000000000000000000000",
INIT_1F => X"8400145AA801741000043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF550",
INIT_20 => X"7FBE8B45AAD568BFFFFAA975FF00003FE0055043FFFFFFFFFDFEFA2D56AB45AA",
INIT_21 => X"F7843FEBA55557FFEFA2D168B55AAFBFFFFFFF80021EF0855421EF00043FFFFF",
INIT_22 => X"A5D2A82155F7AEBFEBAFFD56AA00A2D568B45000002010552EBDF45A28028A00",
INIT_23 => X"BAA2FFC00000804154AA5D00001EFF78428AAA007BC2145F7D5400000004020A",
INIT_24 => X"410AAAEBFF55AAFFC00BAF7AE80010082E954BA0004174AAAA8428B45082ABFE",
INIT_25 => X"0000000000000000000000000000000000000000002E800105D2A95410002A95",
INIT_26 => X"00038F7DB6FBD7490E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA55041549214000",
INIT_27 => X"1F8FD7AAD16FB6DBE8E00155BE8015410140A3FFFFFFFFFDFEFE3F5FAF45AA80",
INIT_28 => X"5B471C7140438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE1049043FFEFE3F",
INIT_29 => X"124BFF7DB68A28A38F7803DE82495B78FC7AAD56FB6DBEF1FAFD7E384001EF14",
INIT_2A => X"FFD1420381C0A02082492A85155E3A4BDE92FFD56FA28B6DF68B551C0E050384",
INIT_2B => X"ABE8E28B7D1420BDEAAA2F1C7038140012482550E021C7EB8028A821C7BC516D",
INIT_2C => X"00492495428082E95400AAA0BDF7DB6F5C70BAFFAE870280024904BA1400174A",
INIT_2D => X"4BA550415410550000000000000000000000000000000000000000000002A850",
INIT_2E => X"DFFFAAD168B55AA80000BAF7FFFDF55002ABFFFFFFFFFFFEFF7FBFDFFFF7AA97",
INIT_2F => X"3DE0000043DFEFA2D56AB45AAD57DFEFF7AA82155F78015400552ABFFEFF7FBF",
INIT_30 => X"568B55A280021EF557FD7555550428B55AAD168B55F7FFFDFEFFFAA955555500",
INIT_31 => X"FBEAB45552E954BA08003DFFFFFAAA8AAAF7843FE10007FEAB55A2D17FFEFFFD",
INIT_32 => X"A842AA00557BD75EFF7D1400AA5D2A82000002A95545A2843FE00F7D17FEAAF7",
INIT_33 => X"0004020AA5D04154BAF7AEA8BEF55003DEAAA2D5554BA5504000105D2A80145A",
INIT_34 => X"0000000000002E974000800154AA002E95410AA843FFFFF7D5554BAF7AE974BA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000002000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000010228001000000000000000000024001620280000000000354200004008",
INIT_04 => X"00016200001310090090004840004152C7208802590000388000004C08006000",
INIT_05 => X"1621008008100002641C0803804000702000000000E02000009900000000B100",
INIT_06 => X"00A0010210200C00000000000000000000000080000000000000D82000000000",
INIT_07 => X"010084C00D267001B880080700285020020AC988200228024004804050089011",
INIT_08 => X"0E0E00000000000000106009872048400C4000010D000008000204150A00815A",
INIT_09 => X"022A040000000000000004C80000002C30C20000000002180800580000000000",
INIT_0A => X"0007600000000000000000080025860000000080A00020602040800000000000",
INIT_0B => X"031400C002000000000000000000000000000000000000000000000000000084",
INIT_0C => X"28DC0D385598035D0008A003B05598035D0008A0034078104B41A41000000000",
INIT_0D => X"041124505598035D0008A000B05598035D0008A0004263C0343EDD4140040422",
INIT_0E => X"B740500401180DE053A98F6ECC739D8140040231068187C39F5A4F985C008902",
INIT_0F => X"000010227848D4303807FC8CC5508AEAED1BFBD406451B02000E033263C0343C",
INIT_10 => X"D6480000000018A700FCF980CC300318A2420851546B2400000040D8549B5800",
INIT_11 => X"81C21140E40511802208D6B30C48F8A8A452210402120A936B0000000004C2A8",
INIT_12 => X"F9E9410006362A2B6424287B08286208D6B1427ED430B41402D0250823597001",
INIT_13 => X"0002C040000000000000000010030060009C000018440021011821B35254E99A",
INIT_14 => X"000040002000044000000000000000000002F0001F00002024B2000200000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"00000000000000000000000000008C8000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C30C30D0A208C4DC822EC1534D34C01FA3F0C7010C6600A0200441920000000",
INIT_1B => X"26130984C26130984C30C30C30D34C30C30C30C30D34C30C30C30C30C30C30C3",
INIT_1C => X"000130984C26130984C26130984C26130984C26130984C26130984C261309A4D",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D00000000000000000000",
INIT_1F => X"AA974BA5D517FFFF08043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA007",
INIT_20 => X"FFFFFFFFF7FBFDF55A28402000F7D56ABFF557BFFFFFFFFFFFFFFFFFBFDFEFFF",
INIT_21 => X"AA8017410007BFFFFFFFFFFFFEFF7D16AB45AA8002000F7D5575455D043FFFFF",
INIT_22 => X"5AAD568B55F7AE955FFAA840201008043FFFFFFFFFDFEFA2D56AB45AA8400145",
INIT_23 => X"FF5D043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE00557BFFFFFFFFBFDF4",
INIT_24 => X"FFFFF80021EF0855421EF002ABFFEFF7D168B55AAD17FFEFF7AE975FF00557FF",
INIT_25 => X"000000000000000000000000000000000000000000557FFEFA2D168B55AAFBFF",
INIT_26 => X"954AA5504154921471FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA55000008255000",
INIT_27 => X"FFFFEFF7FBFAFD7E3A4954BA555B7AFC7080E3FFFFFFFFFFFFFFFFBFDFEFFFAE",
INIT_28 => X"DF52545550A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD74975FFFFFFFF",
INIT_29 => X"AD16FB6DBE8E00155BE8015410147FFFFFFF7FBF8FC7EBD568B55A28000000FF",
INIT_2A => X"497BFDFC7E3F1FAF55A2DB6FB7DF7AE955C7BE800000008043FFEFE3F1F8FD7A",
INIT_2B => X"7EBA0955FF145B7AFC7410438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10",
INIT_2C => X"C7AAD56FB6DBEF1FAFD7E384001EF145B471C71424B8FC7E3D56AB6DB6DF7AFC",
INIT_2D => X"4AA550002000550000000000000000000000000000000000000000000005B78F",
INIT_2E => X"FFEFF7FBFDFFFF7AA974BA55041541055517FFFFFFFFFFFFFFFFFFFFEFF7AA97",
INIT_2F => X"FDF5500517FFFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB45002ABFFFFFFFFF",
INIT_30 => X"56AB55A28002000F7FFC2155552ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FF",
INIT_31 => X"043DFEFA2D56AB45AAD57DFEFF7AA82155F78015400557BFDFEFF7FBEAB55A2D",
INIT_32 => X"FAA9555555003DE00007FFDF45AAD568B45AAFBFFFFFFFAA95545F7840201000",
INIT_33 => X"AAD16ABFFFFFBEAB45A280155EF557FE8B55000428B55AAD168B55F7FFFDFEFF",
INIT_34 => X"0000000000007FEAB55A2D17FFEFFFD568B55A280021EF557FD755555042AB55",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000004000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"0001E6000053300B00D0005800000000000000407B0004BB830004DC3D01E000",
INIT_05 => X"FEE0000008720043EC3C3D0F87FA19F7E0201C409BE1F10623BB000A100CF300",
INIT_06 => X"00200006102FFC8E0007C00078008000171175A200096404D97FFBE4744200AA",
INIT_07 => X"000000482491301000010001DC00000000000000004203FE4005800000008030",
INIT_08 => X"40800020E2008000027FEFF946058180010429000001080AAA010F8000000000",
INIT_09 => X"03EAFE400000120000913FD80000003DF7DE0080010047FBF8000000000800C5",
INIT_0A => X"0800000080000010000400080FFDBE0000004000000100000100506002204610",
INIT_0B => X"FF14FFC00600000000801020000000000000010240001721214E000004000000",
INIT_0C => X"A70C0008020000200000000F30020000200000000F3008001E00000000001803",
INIT_0D => X"004A58F0020000200000000F30020000200000000F3040200000020000000026",
INIT_0E => X"000000000019B140000800800000020000000030B86000400080000200000000",
INIT_0F => X"000014AC08000000508001030A0A4001000000000002183E61E6000040200001",
INIT_10 => X"0000000000A56000090100000000001F86C00010080000000000525801000000",
INIT_11 => X"0600000000001716800000803102020000000002BC360020000000000292C010",
INIT_12 => X"06049CDF70C08040100000706707600000801000000000000057450000100106",
INIT_13 => X"000ADFC011001C81080001101F977FE008000000000000400400400020000805",
INIT_14 => X"0000000000000000000000020020029000000000000000020000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000002000200000000",
INIT_16 => X"0080800801810100000000000093ED8000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000401",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"18618640C49821201C0001A1E79E79A4B0038200010089054C1A0104D2040020",
INIT_1B => X"0C86432190C86432196596596596596596596596596596596596596586186186",
INIT_1C => X"00086432190C86432190C86432190C86432190C86432190C86432190C8643219",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA5504020100800000000000000000000",
INIT_1F => X"AA974AA550002000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7",
INIT_20 => X"FFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFFFFFFFFF7",
INIT_21 => X"5D517FFFF087FFFFFFFFFFFFFFFFFFFFDFEFFFAE974AA5D003FE005D043FFFFF",
INIT_22 => X"FF7FBFDFFFAA84000105D556AB55557BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA",
INIT_23 => X"EF08043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55003FFFFFFFFFFFF",
INIT_24 => X"B45AA8002000F7D5575455D2EBFFFFFFFFFFFEFF7FBEAB55A28000010F7D16AB",
INIT_25 => X"0000000000000000000000000000000000000000007BFFFFFFFFFFFFEFF7D16A",
INIT_26 => X"954BA550000082557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA55040002800000",
INIT_27 => X"FFFFFFFFFFFDFEFF7AE974BA5500050380071FFFFFFFFFFFFFFFFFFFFFFFF7AA",
INIT_28 => X"0038E285D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA55041549214043FFFFFFF",
INIT_29 => X"7FBFAFD7E3A4954BA555B7AFC70871FFFFFFFFFFFFFFF7FBFDFFFFFAA974BA55",
INIT_2A => X"490E3FFFFFFFFFDFEFF7F1FAFC7A28002028555F6FB7D5D75FFFFFFFFFFFFEFF",
INIT_2B => X"5A28402010FFDB6ABEF140A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7",
INIT_2C => X"FFF7FBF8FC7EBD568B55A28000000FFDF525455524BFFFFFFFBFDFC7E3F5E8B4",
INIT_2D => X"4AA5504000BA080000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFEFF7AA974AA550002000557FFFFFFFFFFFFFFFFFFFFFFFFFFAE95",
INIT_2F => X"1541055043FFFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08517FFFFFFFFF",
INIT_30 => X"FFFFEFF7AE974AA550028AAA5D2ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA5504",
INIT_31 => X"517FFFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB4500557FFFFFFFFFDFEFF7F",
INIT_32 => X"A80000BAF7FFFDF55002EBFFFFF7FBFDFEFFFD568B55A284020BA557FFFFFF5D",
INIT_33 => X"F7FBFFF55A2D16AB45AA8402000F7FBEABEF5D2ABFFEFF7FBFDFFFAAD168B55A",
INIT_34 => X"0000000000007BFDFEFF7FBEAB55A2D56AB55A28002000F7FFC215555043DFEF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"1094EC681244819000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"0001E6000053300F01D4587800446194F49020107F0012BBC00202DC3823EA82",
INIT_05 => X"FFF201B228704123FC3C381F87C03DFFF012412A9FE1E01013BF09404050F300",
INIT_06 => X"100B3096F43FFF002004020044041084CB01AD0000037617027FFFE050000080",
INIT_07 => X"A12034043C802A821D41412001A0040950AB60014114C3FE4187A009A663A680",
INIT_08 => X"7F40002C01004000047EFFF811A46968004060629A0002208A00000068113205",
INIT_09 => X"E3EBFE0A812D8D5B742D3FF84056383FF7DE0880042107BFF9C45B85101C49A3",
INIT_0A => X"02804A08221890004806C0310FFDFE00040009814C089202225412115414601D",
INIT_0B => X"FF56FFC0281280080180B2948004400220011100841200D001000624000100C0",
INIT_0C => X"50025360694101816002D41A4068C101815004D8158809C86065941840B1014F",
INIT_0D => X"82418A0068C101816002D41A40694101815004D815810D42E04A08A80098C024",
INIT_0E => X"1A300012682960828F05C96A001B029010134160C8125B0B271802242880A044",
INIT_0F => X"49F115100920C54E8EA256ECF078BA081C10080E05C0B06AA8B12CFD0D42E044",
INIT_10 => X"5144104F30A8801406D00290006280320100010362A8A20826A88660D86B2020",
INIT_11 => X"8010602011819E290048A2118EC8140C08064802C0081B0D64040936443306C5",
INIT_12 => X"C322A4C40A0300600C0A80509F418008804581BA0038005A706680012280506A",
INIT_13 => X"18DBFFC000120080002341881F3FFFF80DCC158092C044600466208CC5091011",
INIT_14 => X"806520398C6021569249C4B3007127080806FF917FC30010107688862A28C545",
INIT_15 => X"9228D9228D9228D9228D9228D99146C9146C84006309044081A001B188300E20",
INIT_16 => X"0448008004000000E07008010003EF80022A51904595123203040D9228D9228D",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_19 => X"0000000000000000004010040100401004010040100401004010040100401004",
INIT_1A => X"7DF7DF7FEFFDFDFFFBE7F3FCF3CF3FFF6EFF7FFDF7FF3EFC1FBFFDF7E0000000",
INIT_1B => X"FEFF7FBFDFEFF7FBFDF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF",
INIT_1C => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFD",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D00020000800000000000000000000",
INIT_1F => X"AE954AA5D00020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"55000200000003FFFFFFFFFFFFFFFFFFFFFFF7AA974BA5D0402000557BFFFFFF",
INIT_22 => X"FFFFFFFFEFF7AE974BA5D00174BA00003FFFFFFFFFFFFFFFFFFFFFFF7AA974AA",
INIT_23 => X"BA5D043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFF",
INIT_24 => X"FEFFFAE974AA5D003FE005D2EBFFFFFFFFFFFFFFFFFFDFEFF7AE954AA5500174",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFD",
INIT_26 => X"974AA550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000001000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"04050005571FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082557BFFFFFFFF",
INIT_29 => X"FFFFDFEFF7AE974BA55000503800003FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D",
INIT_2A => X"140E3FFFFFFFFFFFFFFFFFFDFEFF7AE954BA5D00154AA00043FFFFFFFFFFFFFF",
INIT_2B => X"FFFAA974BA5D00104925D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492",
INIT_2C => X"FFFFFFFFFFFF7FBFDFFFFFAA974BA550038E285D2ABFFFFFFFFFFFFFFFFBFDFE",
INIT_2D => X"4BA5D00000100000000000000000000000000000000000000000000000071FFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02000557BFFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7FFFFFFFFFFF",
INIT_30 => X"BFDFEFF7AE954AA5D041740055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5500",
INIT_31 => X"043FFFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08043FFFFFFFFFFFFFFFF",
INIT_32 => X"7AA974BA550415410552ABFFFFFFFFFFFFFF7FBFDFFFFFAA974AA5D00174BA08",
INIT_33 => X"FFFFFDFEFF7FBFFFFFF7AE954BA5D0000010552ABFFFFFFFFFFFEFF7FBFDFFFF",
INIT_34 => X"000000000000557FFFFFFFFFDFEFF7FFFFFEFF7AE974AA550028AAA5D2EBFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"8632CA211E4491D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"24B000808800040439245B221373581F97B0A8D1040F92000F42000047A00E58",
INIT_05 => X"011B2BBA308F023810004700083E220811E9BF2844021B1004045E4249500449",
INIT_06 => X"EF018980A51003AA0200C020088E16A85235722940A817251100040D6D0702A2",
INIT_07 => X"24E8145C9ECAB0D247B013B405EAD525FAE48FC2060B880081A26DCD4047EFF9",
INIT_08 => X"0050482D0141C0055280100751096B6A40D6F86723E510AA2004803D3275EB20",
INIT_09 => X"20110204804818CD280100207246A8020000AC0283002004051507A5411C0DA0",
INIT_0A => X"4E506A2C6898B2950AA6D635B00041C23020131A80CFDFF3FE509A907C556828",
INIT_0B => X"002200050F60E220A06880D2A14050A028501428054278142151262CA5034385",
INIT_0C => X"F06273612B3482C0C0078E1F412B1582C090078E1F840A2B0114020104022460",
INIT_0D => X"C2C0DB012B1582C0C0078E1F412B3482C090078E1F891C239F8908003099C1AC",
INIT_0E => X"0828041BA859F213AFC14AA380430060181BA1B0FD16770236A4091621C08055",
INIT_0F => X"095337B08AA600CA88B143AB11880C280600101F09C030AB28B03C111C239F87",
INIT_10 => X"3096004B61BD8068B92400D0004E30368910E8822A984B0025B0DE6089462660",
INIT_11 => X"F07830001AC2173B00E162563454C40804055412D4481128C4CC012A66F30455",
INIT_12 => X"BF006850840180A00E1C81900C4190E160589C48082C006A9057CA4385809520",
INIT_13 => X"39C020004416B105036B4180C000800C8C00460848952220592745AC11A544B1",
INIT_14 => X"103D2A512C6A8C4F0008AA800470370000A0004D0000002126F30C902A29C545",
INIT_15 => X"C2A81C2A81C2A81C2A81C2A81C9540E1540E001400006100003202D040050220",
INIT_16 => X"45E22022365034A8EA754008004C0214202C50013456520CA09281C2A81C2A81",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"0040100401004010040100401004010040100401004411044110441104411044",
INIT_19 => X"0000000003FFFFFFFF9004010040100401004010040100401004010040100401",
INIT_1A => X"3CF3CF7FE7FDFD7DF7EFFDDDF7DF7DF7DEFE8FF1F7DEBD6FCD9F7DF7D0512289",
INIT_1B => X"FE7F3F9FCFE7F3F9FCF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"0007F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04000000000000000000000000000",
INIT_1F => X"AE974BA550000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D00020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00000AA007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAA954BA5504000AA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA",
INIT_23 => X"BA5D7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFF",
INIT_24 => X"FFFF7AA974BA5D040200055517FFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500000",
INIT_25 => X"000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040200008000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"00020BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D",
INIT_2A => X"5571FFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5504020AA5D7BFFFFFFFFFFFFFFF",
INIT_2B => X"FF7AA974AA5D00070925D71FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082",
INIT_2C => X"FFFFFFFFFFFFFFFFFFEFF7AA974AA5D040500055517FFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D040200008000000000000000000000000000000000000000000000003FF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAA954AA5D00020AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504",
INIT_31 => X"7BFFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7BFFFFFFFFFFFFFFFFF",
INIT_32 => X"7AA974AA55000200055517FFFFFFFFFFFFFFFFFFFFEFF7AA974BA5504020BA55",
INIT_33 => X"FFFFFFFFFFFFFFDFEFF7AE974AA5D00154105D517FFFFFFFFFFFFFFFFFFFFEFF",
INIT_34 => X"000000000000043FFFFFFFFFFFFFFFFBFDFEFF7AE954AA5D041740055557FFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"5886C0201A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"0005EE040057700F40D08078500000D9218020407F0000BB8018A2FC380BEAC2",
INIT_05 => X"FFE0419028700023FCBC385F87C0BFFFE0124002FFE1E0C517FF09111212F300",
INIT_06 => X"DF0AF116D03FFC96102081020000020489019C4304802412027FFFE000000000",
INIT_07 => X"B710000001160A003475C8100123400E20E1F40F439647FF4807E189A477EF81",
INIT_08 => X"7F0F94801008000007FEFFFB110140695812CC4188D58A0AAA10803448D0844F",
INIT_09 => X"C3EBFD4201258112D4487FF8001010FFF7DE4000000003BFF8C2581808002001",
INIT_0A => X"0801000C024000004A9400000FFDFF50010103134CAFDF03BA18000F39900037",
INIT_0B => X"FF57FFC02812F00429DC92C40002000100008000105400C00400100000A01800",
INIT_0C => X"424202A1CAF13F214001521001CBF03F21100152100801C17E61841950B1C10F",
INIT_0D => X"420B8001CBF03F214001521001CAF13F2110015210088528E00E02C8200A430A",
INIT_0E => X"12480202C86040902AC60BACDF0E02D02001C1C044006D0C94FB94320880603C",
INIT_0F => X"09B00300010AF5052419D196441902801430182800A018D9CA8000648528E00D",
INIT_10 => X"C140004D101808458A5602E000892029110445C19960A00026880C0067390000",
INIT_11 => X"4040301009408021144CB042F880100C0601844068880CE72000013600600332",
INIT_12 => X"EE38A1F80E02120018390320F050144CB241D0B9023402085020825132C8CB5B",
INIT_13 => X"001BFFC200400020224000405F7FFFE0008E17C0D240406519400500840A9524",
INIT_14 => X"907120AC810033149249C433200180082A06FF907FC308181204800600000000",
INIT_15 => X"1010C1010C1010C1010C1010C10086080860840063090442A18001B188300C48",
INIT_16 => X"2000100100000000000004002403EFC10302219A41C1443243050C1010C1010C",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_19 => X"0000000000000000000080200802008020080200802008020080200802008020",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"550000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974AA550400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"00087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE954AA5D00000AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA5504020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA55",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400010087FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE954AA5D0402038007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE954AA5D00020BA087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"00010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D00",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA55040001000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAA954AA5D04000AA087FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D00020AA007BFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"0000745C200801000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"0001E6000053300F00D0007810042140C00000407F0000BB800000DC3801EA00",
INIT_05 => X"FFE0000008700003FC3C380F87C019FFE01240009BE1E00003BF00000000F300",
INIT_06 => X"DC8C3006103FFC0000000000000000048900880100800012027FFFE000000000",
INIT_07 => X"0061200009B24B043980021000810284204A8001401643FE4007E5501AA00000",
INIT_08 => X"7F00000000000000007EFFFB11A56940581280031D61420000B080102040BC5B",
INIT_09 => X"C3EBFC020125811254083FF80000003FF7DE0000000003BFF800580000000001",
INIT_0A => X"0580000000000000000000000FFDFF4000000AA0354000019C40000128000011",
INIT_0B => X"FF56FFC000104000000010440000000000000000001000C00000000000000240",
INIT_0C => X"48C0804012500021B00880108012500021E00880104809C1666594584031010F",
INIT_0D => X"0501840012500021B00880108012500021E0088010492064206100E810842000",
INIT_0E => X"0270040410004C840041A0D8005410903804100144800803419043064900C002",
INIT_0F => X"400041020902F60002260D65B361BAA1041018140F02C0000809408D20642053",
INIT_10 => X"D0021800020818B06D9802F00030C02060110002C9E8010C00010480B35A0300",
INIT_11 => X"90203020042108603100061516EE800C060228204300166B4060080008240593",
INIT_12 => X"14AE4C7C02000040206602C10B48110006143B62023C00142800B04400095DFF",
INIT_13 => X"001BFFC000000000000000001F17FFE000DC1180C78044000440292083010402",
INIT_14 => X"814080008000010012414433000100080806FD107FC300000000000600000000",
INIT_15 => X"1000C1000C1000C1000C1000C100060800608400630104408180012188300C00",
INIT_16 => X"0000000000000000000000000003EF80020201904181003003000C1000C1000C",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"3DF3DF64C7986120B42BB99575D75FFD2AF6E7CC1132CD73DF3A441990000000",
INIT_1B => X"1E0F0783C1E0F0783DF7DF7DF7CF3CF3CF3CF3CF3DF7DF7DF7DF7DF7DF3DF3DF",
INIT_1C => X"0000F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100800000000000000000000",
INIT_1F => X"AE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"00007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D00020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010080000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000001008",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA550000010087FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002010087FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00004000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"4909E6093253306F82D0007C80000000080E01007F8020BBC00040DC3801EA00",
INIT_05 => X"FFE0000008704503FE3C380F87C019FFF01241009BE1E00203BF80800000F392",
INIT_06 => X"CC083006103FFF9E2086C2086E006604C9019D03108B7412027FFFE070400880",
INIT_07 => X"0000004024057000000100000000000000000001401643FE4007C00000000000",
INIT_08 => X"7F00000801404000007EFFFF40010000401408000045000000A0801000408000",
INIT_09 => X"C3EBFF4A7DF795965C6D3FFC0020003FF7DF01880C618FBFFDD75E0010004043",
INIT_0A => X"0000000000000000009400000FFDFFC006020000000000019804000028000191",
INIT_0B => X"FF56FFC02812E0182000F2C48304418220C11160845004D04820000000000000",
INIT_0C => X"0800800002400001000800000002400001000800000801C0786184185031810F",
INIT_0D => X"0400000002400001000800000002400001000800000000202000000800000000",
INIT_0E => X"0200000000000404000000880000001000000001000000000090000008000000",
INIT_0F => X"000040000100C600800001040000040009100000000200200000400000202000",
INIT_10 => X"4000000002000000081001000000000040010000082000000001000001080000",
INIT_11 => X"0000400080000040010000001080001008000000010000210000000008000010",
INIT_12 => X"0420000000030280000000010000010000001020000000000000100400000108",
INIT_13 => X"001BFFE0120012C1400080291F17FFF0018C11808200400000400000C2000000",
INIT_14 => X"80400000800001001243443B000100880806FD107FC301800000000600000000",
INIT_15 => X"1000C1000C1000C1000C1000C10006080060840077330C4889CC292588300C00",
INIT_16 => X"44C82082068C0200000008014023EF80020201904189003003000C1000C1000C",
INIT_17 => X"4110441104411044110441104411044110441104411044110441104411044510",
INIT_18 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_19 => X"2FFFFFFFFFFFFFFFFFC110441104411044110441104411044110441104411044",
INIT_1A => X"0924821409005312E8A25E15A69A6BFB0A196A8C5A2932F7C13C15DA08080000",
INIT_1B => X"C46231188C462311892492492492492492492492482082082082082082092482",
INIT_1C => X"00162B158AC562B158AC562B158AC562B158AC562B158AC562B158AC562B1188",
INIT_1D => X"0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"00087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04000",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040200000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"94A7B2B1450000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"6FEBEF5FEC737AFBC6F85FDEB220109E1FEFFFE3FBA7FDFB9BD301DC3FF5F0D2",
INIT_05 => X"FEEDBFDC387F987FEF7C3FAF87FF59F7F5FB7FF59BE1FF980BBBB7FE6D21F3DB",
INIT_06 => X"DFA08957902FFDEE9D7DC9D7DF2B263893479DDFAFDFE15213FFFBE1F1D3A333",
INIT_07 => X"00018010992310605CE10301DE0C1831CB7DF60A244B9BFEE00589DDBCEFEDC1",
INIT_08 => X"FFEFAA001D8EA111DA7FEFF90F21C8C84D9C0D858FC7020828C18FD18346BBF0",
INIT_09 => X"0BFAFFF37DF7B9DF7DCB3FDE89ECC07DF7DF5F985C6BCFFBFA28F99E7EB07F47",
INIT_0A => X"0607307DCFE1D4077B4D0026FFFFBE7D67D7F3BB79CFFB83BF14EC1E7D598058",
INIT_0B => X"FFFCFFC7D7D51D6F5FDCB935D7AFEBD7F5EBFBF7FEBD66DBFCA3F87501AE7B08",
INIT_0C => X"40520201F45EC0010007E01001F45EC0010007E010084BCD7FF1B61B5C33813F",
INIT_0D => X"0001A001F45EC0010007E01001F45EC0010007E01001BD8020500008001F0100",
INIT_0E => X"0200001EC00040B02007EC09A0E00010001DC0004600400F781429C008000077",
INIT_0F => X"81C203404B3BFD0402346235408402C08010003C064000E408010081BD802060",
INIT_10 => X"68B1000E401A08FE0012040000FC002001360403E434588007200D00F88C84C0",
INIT_11 => X"281D00001F01002156040675809145400007B00040091F1190982038406807C8",
INIT_12 => X"903A80008320C0403C34000088601604067D00212000007C400082D81009FC08",
INIT_13 => X"D6BFDFF7BFFED3FBFF6A84383F177FF005FFBFF5FA1040076065F730FC08043A",
INIT_14 => X"CDEBCFF589807B7096CD4CF73AC1FC98884FFF19FFC71FEFED7B251E35768E8E",
INIT_15 => X"78C0D78C0D78C0D78C0D78C0D7A606BC606B8C56F7730ECCDBDF152199F51EDD",
INIT_16 => X"FEFDFDDFE7DD87FEFF7FF796FFFFFDFFD7E681B867D3683A03A40F78C0D78C0D",
INIT_17 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFB",
INIT_18 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_19 => X"6FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_1A => X"4C30C375E2BD54D5D6C565F871C71D44FCF491E166CC853E8695F86EDB5C8864",
INIT_1B => X"26130984C26130984C30C30C30C30C30C30C30C30C30C30C30C30C30C30D34D3",
INIT_1C => X"000130984C26130984C26130984C26130984C26130984C26130984C26130984C",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"1085B0B041000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"6FAB975B6470BAF386C87A9CB00000001FEF9F23E3A7BDE79B5101D23FB5C0C2",
INIT_05 => X"F8EDBFD4347F18778E723F2E47FE59C7F5FB7F759B91FB880BA3B6FE2921CBDB",
INIT_06 => X"DFC00147000FFC128D5CE8D5CC210638A046889CAB57E84217FFE3E181932377",
INIT_07 => X"000141000000042000000288020C18300320620A80231BFE200181092CE7ED80",
INIT_08 => X"FEEF22000C562551D87E8FF90041101042110180004102800008801183468180",
INIT_09 => X"0BE0FC137FF7A0FF75813F1C85244071EFBF17D85C738BE3FA08F9DE36B05B07",
INIT_0A => X"040510768EA0C406630D00226FFE3E2D62D6E21259CFDB039E806C0245188040",
INIT_0B => X"FF48FFCC57550D63564D1D2556ADAB56D5AB6AD7EAB962CBD8A3A83101F47E08",
INIT_0C => X"00130201E44A40010007600005E44A4001000760000843C561E5C55C42B9011F",
INIT_0D => X"00002005E44A40010007600005E44A40010007600004BD8020100008001F0100",
INIT_0E => X"0200001EC00000382006EC0820A00010001DC0000208400D781020C008000077",
INIT_0F => X"81C20040431BC50402146235400400408010003C064000C400018080BD802020",
INIT_10 => X"4821000E400204FE0010040000FC0000003E0403A424108007200102E8888080",
INIT_11 => X"080500001F0100005E040475808101400007B00000015D111010203840081748",
INIT_12 => X"903A8000012040403C34000080201E04047D00202000007C400000F81001FC08",
INIT_13 => X"109E1FE5ADA4C25ADE72041A3F147FF0018DBBB5FA10400360649310FC08003A",
INIT_14 => X"EFABC7054880693016DD4C755AC16C1A884FFE18FFD757E7ED7A211E81C09818",
INIT_15 => X"3440C3440C3440C3440C3440C3C2061A2061AD46FF730E5CCBCD55219AB55F0D",
INIT_16 => X"DE75ED5EC71385FC2512E3565BBBF1BAD6F281BC63F1683803C00E3440C3440C",
INIT_17 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6B",
INIT_18 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_19 => X"7FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_1A => X"0000003C010072F24388521000000140A8100481CA8604368714104A47168874",
INIT_1B => X"8040201008040201000000000000000000000000000000000000000010400000",
INIT_1C => X"00140A05028140A05028140A05028140A05028140A05028140A05028140A0100",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"8C2100804900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"02000100440408002408008002221000204116A280000F000001400000100010",
INIT_05 => X"0004D44400004D4400000000000000000000005C0000000A0000002C20600000",
INIT_06 => X"2000004100000120040A0040A00B009000620294010000400080000888800911",
INIT_07 => X"2488045002489020420110800244891211440804000810002000081040000000",
INIT_08 => X"00B062080542C004CA00000050080202008401842004108AAAA00008912240A1",
INIT_09 => X"2800010000000C0000E400002040500000009202C10020400044000222000204",
INIT_0A => X"02043058C460540329810002D002000400407020800000004000640800088008",
INIT_0B => X"0008000140000401028008330000800040002002480102010082981500062108",
INIT_0C => X"00500000040A40000000A00000040A40000000A0000040060084104110828030",
INIT_0D => X"00012000040A40000000A00000040A40000000A0000000800010000000000000",
INIT_0E => X"00000000000000A00000040020A000000000000006000000080020C000000000",
INIT_0F => X"8000024040152000000020000004004080000000000000240000000000800020",
INIT_10 => X"0821000000120002000004000000000001220000040410800000090000808080",
INIT_11 => X"0805000000000001420000200001014000000000000900101010200000480008",
INIT_12 => X"0000000001204000000000000820020000200000200000000000028800002000",
INIT_13 => X"29400000933050080C0001900020000000408010000000022000D61028000008",
INIT_14 => X"440245400082D022040000400800081022C0000080000206CB0821082B694D4D",
INIT_15 => X"605016050160501605016050160280B0280B0012000843066021001400040024",
INIT_16 => X"0810840861CD33548542A10209D4100E4040A00002002C004001036050160501",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008021",
INIT_18 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_19 => X"0000000000000000000020080200802008020080200802008020080200802008",
INIT_1A => X"41041001A835050788440B58C30C31DF6C110A00246972C0C39989A40A0C22E1",
INIT_1B => X"C06030180C060301810410410410410410410410410410410410410410410410",
INIT_1C => X"00160B0582C160B0582C160B0582C160B0582C160B0582C160B0582C160B0180",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0803B2814D0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"26E1E905CC574828C4F85FC600000016004F77E2F887CDB80BC340DC07D1F000",
INIT_05 => X"FE1DFE4C080F884FE33C078F803F19F011E93ED49BE01F1A03B8972E6D20F049",
INIT_06 => X"64A08857902000DE142D4142D5030010134395D70589415002FFF800F0C38111",
INIT_07 => X"00088400092300601CE00101DE040811D919F402244293FEE00400CCB46BA4C1",
INIT_08 => X"7FA0AA08148A4000887FE0000F20C8C80D080D818FC2000000418FD08142BAD0",
INIT_09 => X"0BFA02E204D2154D28AA3FC60888D03C10415A80402847F8002458926A002E45",
INIT_0A => X"0406305587A1540231410006DFFF80540541619968C76980E914E4163D498010",
INIT_0B => X"FFFC0007C7C0140D0B50A8218102C0816040B1225C1506512C83E85500AC3A08",
INIT_0C => X"40520000141EC0000000A01000141EC0000000A01008480D3EB4A24A0C910037",
INIT_0D => X"0001A000141EC0000000A01000141EC0000000A0100100800050000000000000",
INIT_0E => X"00000000000040B000010401A0E000000000000046000002080429C000000000",
INIT_0F => X"80000340483B590000202000008402C080000000000000240801000100800060",
INIT_10 => X"28B10000001A08020002040000000020013600004414588000000D00108484C0",
INIT_11 => X"281D000000000021560002200011454000000000400902109098200000680088",
INIT_12 => X"000000008320C00000000000086016000220000120000000000082D800082000",
INIT_13 => X"D6ABC032936E43A92F2880B01F37001004B29450580000066021F6303C000408",
INIT_14 => X"45624DB481806A62840800C22800B8900042FF0180000ABFEF89250815568A8A",
INIT_15 => X"68D0068D0068D0068D0068D006A68034680300021410028450530014014002D4",
INIT_16 => X"2C989489418D13FE7F3FFD8BADB7FC4F4164A00806522C0A40A50268D0068D00",
INIT_17 => X"C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C4B1",
INIT_18 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_19 => X"2FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_1A => X"5D75D7FFEFFDF9FAF3E7E3EFFFFFFEBFD6EE7FFDF7FE78FC3CEFFDFFEA0C0060",
INIT_1B => X"EFF7FBFDFEFF7FBFDF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DD75D75D7",
INIT_1C => X"001F7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDF",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"3CF3CF75EFBD75F5FFEFFDFDF7DF7FFFFEFF9FE1F7FFBFEFDFBBFDFFD0000000",
INIT_1B => X"FE7F3F9FCFE7F3F9FCF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"0007F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"1084B030000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"6DA986092050306382C05A1C900000001FAE89016387B2A38B5000D03FA1C0C2",
INIT_05 => X"F8F92B90307F41338E303F0E07FE19C7F1FB7F289B81FB8003A396D20940C3DB",
INIT_06 => X"DF800106000FFC020004C0004C0006288004880800036002137FE3E101030222",
INIT_07 => X"000100000000000000000220000810200220620E00030BFE000181092CE7ED80",
INIT_08 => X"7E4F400000000001107E8FF90001000040100000004102200000801102448100",
INIT_09 => X"23E0FC027DF780DF74013F1C00240071E79F05888C618BA3F800599C10104903",
INIT_0A => X"040100240A808004420400202FFC3E002202021259CFDB039E00080245100000",
INIT_0B => X"FF40FFC407500020004C10060204010200810040801060C04821202001A05A00",
INIT_0C => X"00020201E04000010007400001E0400001000740000803C0616184184031010F",
INIT_0D => X"00000001E04000010007400001E04000010007400000BD0020000008001F0100",
INIT_0E => X"0200001EC00000102006E80800000010001DC0000000400D7010000008000077",
INIT_0F => X"01C200000308C50402144235400000000010003C064000C000010080BD002000",
INIT_10 => X"4000000E400000FC0010000000FC000000140403A020000007200000E8080000",
INIT_11 => X"000000001F01000014040455808000000007B00000001D010000003840000740",
INIT_12 => X"903A8000000000403C34000080001404045D00200000007C400000501001DC08",
INIT_13 => X"001A1FE004048240426200081F147FF0018C1380DA10400140640100D4080032",
INIT_14 => X"812982050800A91012494C31004124080886FE187FC301B124F2001600000000",
INIT_15 => X"1000C1000C1000C1000C1000C18006080060840477330C4889CC012188310E08",
INIT_16 => X"44602002061004A820104809402BE1900222019861D1403803800C1000C1000C",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"2FFFFFFFFFFFFFFFFF8100401004010040100401004010040100401004010040",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000100080",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"88280C4C7B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"00160090920C04800904848262220277E05152B280780D407428E723C01E1400",
INIT_05 => X"0006D46207801E400183C0707800E6000E008057641E00473C40680D32330C00",
INIT_06 => X"203F70C165000225E2C11E2C12A0D0144AC27206582C166504800000B0FC21D5",
INIT_07 => X"920CFC5E6D233B964E7CD99DFB870E1DDDD889C5FBDC440129A0604442180238",
INIT_08 => X"80B036AD23C17544C581000657A0E8E83D86F0E4A7B2D88AAAFD7FE0E1833AC5",
INIT_09 => X"C800016D82082E2081B6C0027ADA398000008A504318404005B70663212C04A0",
INIT_0A => X"4AF4AA414568729139FAD610C00001A2502440888420247041E87681008CE9AF",
INIT_0B => X"00890022B826E250B12346F1244812240912048941621804A150CA1CA45C254D",
INIT_0C => X"B2E0F1F80FA97FE0F0009E0FC40FA97FE0F0009E0FC048211E9C11C31F82E4A0",
INIT_0D => X"C3CB5F040FAB3FE0F0009E0FC40FAB3FE0F0009E0FCC42EFDFBF0AE03080E2AE",
INIT_0E => X"187806013879BA878FE807F65FBF12E0380231F0BD9E3FC08FEBD6F661C0E008",
INIT_0F => X"C83136B248831ACBFC8BBDCAB779BC699F20180309A0F83BE2B87C7C42EFDFBF",
INIT_10 => X"9947184131B59003FFEC07F00003F01FB90BE9F01FC8B38C2098DAE007F323A0",
INIT_11 => X"D065703080E29F1B2BE9F8A27E6E915C0E004C72BEC800FE7464290626D7003F",
INIT_12 => X"6F846DFC0C2352A0024B83F07F198BE9F8A0FFDA2A3C0202B8776A2FA7F023F7",
INIT_13 => X"11800014481A6105810941C5C068000CD4004C0905E52630BB1AE49C2BA7F98D",
INIT_14 => X"7E96656074EA560F0416A24844B01302A26100C4801844069B0C88881A28C141",
INIT_15 => X"E2781EA781E2781EA781E2781C33C0613C0E21020800239450116ED443C041B4",
INIT_16 => X"8112C1241140A056954AB0C280D0002020187007122C3E04E03383E2781EA781",
INIT_17 => X"1204812048120481204812048120481204812048120481204812048120481205",
INIT_18 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_19 => X"4000000000000000001204812048120481204812048120481204812048120481",
INIT_1A => X"10410411062084E57CE2641DC71C71574E09B56C74DAB16782171CF13043A85D",
INIT_1B => X"F87C3E1F0F87C3E1F04104104104104104104104104104104104104104104104",
INIT_1C => X"0007C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0",
INIT_1D => X"0000000000000000000000000187C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE500",
INIT_1E => X"BD54BAF7FFD55EF007FD75EFFFAE97555557BD75EF5D00000000000000000000",
INIT_1F => X"FFC0000AA843FE00AAFBE8B45AA803DFEFA28428B455D0017410A28428AAAA2F",
INIT_20 => X"57FFFEBAA2D5401450051401555D7FC0145F7AEBFFFF08002AA10A2AABFEAAA2",
INIT_21 => X"5D7BD755555517FFEFA280021FF082E974AA5D7BFFE000804000BAAAAAAAB455",
INIT_22 => X"A5D2EA8B45005168A10AA8028A10087FD7410557FC21555D51574AAA2FFE8B45",
INIT_23 => X"FFFFAE95410AA80000005D003FEAAFFAEBFE00A2803FEBA002A820AA0800174B",
INIT_24 => X"5EFA2AEA8A10000417410A2FFE8BEFF7FFE8B45FFFBC00005D003FF45557FC01",
INIT_25 => X"000000000000000000000000000000000000000000557DF5500003DFEFFF8417",
INIT_26 => X"12555F524AFE38B780154BAFFF1D54AF0075D75EFEBAE9554540754717F1F800",
INIT_27 => X"B6AB50B6AABDE12BEA0AF010B7D1F8F47E00A2DB45AA8A3AFD7B68E2AB78550E",
INIT_28 => X"A43FE9257F1E816D557095EAAA2D1401D500002A150038038E285D7F78FD7000",
INIT_29 => X"57545A87AAD178A8002D1D21C5E8257D5C7AA854008700249243A412EBFF5542",
INIT_2A => X"02D152A82000E3A5D2150AB8F401471EDBC0B680900AAF52B474385D75C502D1",
INIT_2B => X"D417FD7E9541242FE920AD082E10A28F6A150012A2F02AFFDF40E85F475451D5",
INIT_2C => X"55080550E87B7A405B52AAD152BD00151EAFEDB52E3F1EFFFF485A2DA3D5D24B",
INIT_2D => X"445057F40545850000000000000000000000000000000000000000000005AAF5",
INIT_2E => X"AB55F7AEAABFF5D2A81151FB8635A02FA69574BAF7D5555AF0D79D55FFA2AC97",
INIT_2F => X"34A08D46F6ABE7082AAAAF2FAC77FE00FF16565B2FA9075F4F7B3EBDF50FEAEA",
INIT_30 => X"C95256803CE3AEB038662E5D81406014D5D51F5E08A394003A908B8410E707EF",
INIT_31 => X"C0954AF0151555AF58794040077D774FAE8C798A11A0EAEF75F7AA84001A7052",
INIT_32 => X"245B4E1870108B11020AD4AA05542A0A05051023F9A9D57B63BFBF906CB45FAB",
INIT_33 => X"ABD5F5F0DA6BC9525688C1A2A0C06E9FEE5555BE48AB2A2AE0A0F20C43EAC562",
INIT_34 => X"0FF8000000FF80F55E25C00A0BA7FBED407A97F6F35F498B96BEB12DAAB77558",
INIT_35 => X"00FF8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF800000",
INIT_36 => X"000000000000000000000000000000FF8000000FF8000000FF8000000FF80000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000800000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"CA1800080848B0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000010822C00803804000001999EF9C00040B0002000001000640200001018",
INIT_05 => X"0000400244000000014200004000000004000000001000032000200002100800",
INIT_06 => X"202800208500000080412804100CB08000302220080408010000000404100844",
INIT_07 => X"25FC4C5AF6FEF002230018010860C1833C460044204C000008A0041000080008",
INIT_08 => X"0010008D22C0F55000010000524481890BC000263000188AAAA10F8C1830562B",
INIT_09 => X"041001B102002E20013600022D8819000000A000110A4000002C204000240420",
INIT_0A => X"0BE0B002605C1C1108484400C000002040040820000020104100028800002801",
INIT_0B => X"000000081001004010810510040802040102008100200800A1100707040101E2",
INIT_0C => X"10F18058000003C0F000A000C4000003C0F000A000C0000012187087010AE4B0",
INIT_0D => X"00012704000003C0F000A000C4000003C0F000A000CC4200002F08E030800000",
INIT_0E => X"1878060000000AAC00680000001F10E038000000078808C00000023461C0E000",
INIT_0F => X"4800025200040A00D000000202090C281F201803000000240218C0044200001E",
INIT_10 => X"904618400012900001EC03F000000000392100B00048230C200009A000130320",
INIT_11 => X"806070308000000961002880204A901C0E00000002C9000260640900004D0000",
INIT_12 => X"0904285C0C0312A002000000083881002880025A0A3C020000002A8400B00007",
INIT_13 => X"08400004080030008010468220A00008D0000801046004308A18500002012800",
INIT_14 => X"2200000840280206089000004090110200000000001454000200828008081110",
INIT_15 => X"A4191A4191AC191AC191A4191A00C8560C8D2910000060901010401E13405111",
INIT_16 => X"8000410410028000100800140000002004103224002006406401918C191AC191",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"0000000000000000000200802008020080200802008020080200802008020080",
INIT_1A => X"1451455901218D2C4CA2900C9249258306BABEFC54A081701C397452B4008A04",
INIT_1B => X"BADD6EB75BADD6EB755555555555555555555555555555555555555545145145",
INIT_1C => X"0005D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2EB75",
INIT_1D => X"0000000000000000000000000607FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF600",
INIT_1E => X"E80010AAAABFFFFFF803FE10F7D17FEBA55556AAAAAA80000000000000000000",
INIT_1F => X"2EBFEBAFFD555400557BD54BA5D7FFDF45A2FBD75EFA2AE97555F7FBFFF45FFA",
INIT_20 => X"A802ABEFA2D568A005D5157400AA8028AAAF7FBD54AA002A955555D7FE8ABA08",
INIT_21 => X"FFFFFDF55AAFBC0010555540010550417555AA8028BEFAAAE97555082A80000A",
INIT_22 => X"A557BD7410550428ABA5D5168ABA552EBDFEF5D7FEAA00AAAABFEAA007BC0145",
INIT_23 => X"FFFFFFEAB55557FFFEBAAAD568B45A2D5575555D7FC2155F7AEA8BEFAAAA954B",
INIT_24 => X"4AA5D7BD74000804154BA082ABFF55FFD57DF45F7D568ABAF7AABFFFF082ABFF",
INIT_25 => X"0000000000000000000000000000000000000000002EBFFEFA280021FF082E97",
INIT_26 => X"95545E175EFF57BF8FC2000BEA4BAE97F78A3FE28E3D17DEAA485FE8E02B5000",
INIT_27 => X"FD55455571E8A2A087BF8EAAEB8E0016D5D75D54BA5D7BFFF7DA2FFD55EFAAA4",
INIT_28 => X"AA07157428145A00AA8A2FBD7B6DF6AA28550E10405F7A4AFE38EAA0924921C2",
INIT_29 => X"6AAB8E971471C7010B7D168F47400A07A28415A001684104155C5B6DF6DBEFBF",
INIT_2A => X"5FD4BFBD7B6A0BF492415FC20105D24AAABF1FFBC7010FF8A38FEF557FEAB78B",
INIT_2B => X"FE38017EBA4A8EB8F6FFD5FE8B7D557495EAAA2D16D1FDBED56A55557A43DE38",
INIT_2C => X"C7AA854008700249243A417FFF41542F5D717FE2AAAA56DEBD17FE3DF7FB7FEB",
INIT_2D => X"FBA007DFCA127B8000000000000000000000000000000000000000000002A3D5",
INIT_2E => X"FFEFAAFBD55FFAA8416545A6FB60F47AF2A00010F78028B15F7823FEAAA2D57D",
INIT_2F => X"21A022A38C20B2552E975F758516AAAA0869AAAB8A7C19C55550E8574BA557BF",
INIT_30 => X"895755FFEFBCEE5FBAACB10085EE5DE10A2AEBFF55F7BAAA8565DBAC1112FFAC",
INIT_31 => X"02EABEA097BEAAFAF2863FA00DD574201E7AD1FFF5575841DE08007FC2048002",
INIT_32 => X"AF9554FF57EFBFA18D4FBFFF40FF809D4000D7FC00FC5D062BBA05ED5034472A",
INIT_33 => X"FED17DFBFF6963FCAAA2283CF14050062B0A2F7AE8B5D5D51F5E18ABD5EAFFF2",
INIT_34 => X"0000000000002CB75F7AA84001A7052C95256807DC31AA8114DE55F5BED201FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000800000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2812",
INIT_01 => X"0005A18A0849204D1CA024A542500368404000720885800802000106E4D10204",
INIT_02 => X"5C010802020408040C600850AA055254090541A111240A104A0000000908B510",
INIT_03 => X"182202210800004401060A0010041028021560A0218808002440840008C80550",
INIT_04 => X"21030A008814500120A06B0870201010258261E141A2326511024182142494D2",
INIT_05 => X"48484098142953388552102442884882B58A09291290A1120A81A3C200418DCA",
INIT_06 => X"22208802800554529001C9003A2800203120000104810100002A614008102244",
INIT_07 => X"0008040000221040408100890C0000011804480420420154000088096A0EA8C0",
INIT_08 => X"B846C0081190C105424705510A08828A0B190C0428040080A0A10F8000009200",
INIT_09 => X"20B0573165541CD54822160A89E89020AA8A80CA9D39CE215264B15818004442",
INIT_0A => X"0402100C088104010AC80005C568147007031012D40D71824114081538000048",
INIT_0B => X"550055481205100C000134128304408020C11020040244D00001306100A24600",
INIT_0C => X"00500000B01480010000A00001501480010000A0000801487334E34C1A980001",
INIT_0D => X"00012001501480010000A00000B01480010000A0000138000040000800000000",
INIT_0E => X"02000000000000A00003600180400010000000000608000A5004090008000000",
INIT_0F => X"000002400008C4000220420040800280001000000000002400000001A1000040",
INIT_10 => X"2090000000120C94000200000000000001380001C01048000000090298040440",
INIT_11 => X"2018000000000001580002508010440000000000000953008088000000481380",
INIT_12 => X"10180000820080000000000008201800024C000100000000000002E000095000",
INIT_13 => X"09130A82000C90A0000081A004342AB001720040000000000001502050000422",
INIT_14 => X"094882958000934200904407600090822085E0100D52498002B1041092001514",
INIT_15 => X"3C1011C1013C1011C10134101140801A0808AD4451394CD0391A541593C04B59",
INIT_16 => X"022810800000A0289A6D084D4021208106142034406144004041011410114101",
INIT_17 => X"4010040104411044110441100401004010040104411044110441100401004010",
INIT_18 => X"0102401024010241106411064110640102401024010441104411044110040100",
INIT_19 => X"2F81F81F83F03F03F04110641106411064010240102401024110641106411064",
INIT_1A => X"0820823047486021658010816596597700138D70C030B542923650C7D0002281",
INIT_1B => X"944A25128944A251282082082082082082082082082082082082082082082082",
INIT_1C => X"F804A25128944A25128944A25128944A25128944A25128944A25128944A25128",
INIT_1D => X"0000000000000000000000000787C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF871",
INIT_1E => X"5420AAAA843DFFFAAD1554005D7FD74AA0004001550000000000000000000000",
INIT_1F => X"2EBFF45AAAAA8A10A2AE80010A2AA975FF5D003FE10F7D17FEBAF7D5420AA085",
INIT_20 => X"D7FFFF45A2AA975EFA2FFD7555FFFBFFF45AAFBC20AAF7D1575EF55517DF555D",
INIT_21 => X"AAAE95555552E974105D517DF55AAAAAABEFAAD1575EFAAAE974AA5D51554BA5",
INIT_22 => X"F552E82010F7AABFE10FFD542145FFD5554AA555555555557FE8ABA082EBFFFF",
INIT_23 => X"EFF7FBC0010AA802ABEFAAD540000FFD540000AA802AABAF7FFC2010AAAE821E",
INIT_24 => X"555AA8028BEFAAAE821550851420AA002E800AA08042AB45007FC00BAFFD168B",
INIT_25 => X"0000000000000000000000000000000000000000002E80010555540010550417",
INIT_26 => X"7DEAAE95F40002157F470AABE803AE97A2DF55400557FD54AA1D04001C515000",
INIT_27 => X"E105EF55517DFC5552ABDF45B6AEAFFD5F7A482000BEAE905C755003FE28E3D1",
INIT_28 => X"A4070BA5FD0154BA5D7BFAF7DA2AE955EFAAA495545E3F5EFF57F7FE80082FFD",
INIT_29 => X"571E8AAF082AB8EAAEB8E0016D5D2A924105D5B7FF7DB6AAAABC7BEDB505EFBE",
INIT_2A => X"E80495038AAAEAF1D7410E80000FF8438E00B6DF68FEF4871D24BA495B5556D5",
INIT_2B => X"80071ED1EFEAF1EFFFDEAD1C5010AA8E2FBD7B6DF47A00EBDB50000A380AAE28",
INIT_2C => X"28415A001684104155C5B68E2DBEFBFFBC703AE2DF42AAA002A851C214003FF6",
INIT_2D => X"4AA550002155510000000000000000000000000000000000000000000002087A",
INIT_2E => X"215555003FEAAAAD57DEBAA2FDDC01051FBD74BAF7802AB05AAFBD5400557BD5",
INIT_2F => X"60F47AF7FC20B2F7FBC015D58517FF555D2ABDF55F782BEB47AFAD00010F7AA8",
INIT_30 => X"22A955FFFFC20FFF3AE544108410174BA557BEABEFAAEBD55FFAA1456547A2D3",
INIT_31 => X"D4420BA547FD75FF58516AAAA0828AAAB4A78016545540400010557BFDFFFF78",
INIT_32 => X"FFBD550AAFACAAA122AA8954BAA2AE9D545002A800A8FF862BA00F2F9E8F0050",
INIT_33 => X"002E954505C417FFFF08555555BAAD335B57AB5155400A2AEBFF45FFFB404007",
INIT_34 => X"000000000000061DE08007FC2048002895755FFAEBCFE57BBA57002DF3C4AAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000001000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B815602110494074133520400E02B92206",
INIT_01 => X"014C9BC048800168240442C99E004B61404040028804A0080A000516A0990A08",
INIT_02 => X"4809A900031800444440589866E331352180D468B8000E600C0081110B802CD0",
INIT_03 => X"DA16C0200C0001423583480408D60520320066810A80881068A808029C856330",
INIT_04 => X"2088681DA82740EC92307364B37569100A84E1E11C251210990040420E005A48",
INIT_05 => X"2D284A102414411A314A0A02C18C01B9854368280A506902018C2442484038D1",
INIT_06 => X"23600016801CCCAA9061C9061C0D0080001005210C8761001166CCC40C110826",
INIT_07 => X"0178045800B6540063000889082040A13A0716042440833280038C89904E6400",
INIT_08 => X"D20A480810804451421D1CC8024481994B5500061000088000A10F840854973A",
INIT_09 => X"2079CCB035E03CCC5D2A35620988100A698761C0953B6E84C82C404018304D42",
INIT_0A => X"070070202A90340440C80004CCE4CC1042061913208CE8024380880820010040",
INIT_0B => X"3302CCC01300104018900402870C4287214210E114200410EC20242D01015E84",
INIT_0C => X"4801000180148000000800100040148000000800100401C33249049051218073",
INIT_0D => X"04008001001480000008001000E014800000080010001C000040000000000000",
INIT_0E => X"0000000000004408000068018040000000000001400800091004090000000000",
INIT_0F => X"00004100812644000004400140800280000000000002000008008000B0000040",
INIT_10 => X"20900000020800CC0002000000000020400800030010480000010400C8040440",
INIT_11 => X"2018000000000060080004418010440000000000410015008088000008200540",
INIT_12 => X"80188000820080000000000100400800041C0001000000000000902000014C00",
INIT_13 => X"284B264208448260E27285A23224E660084208410000004444000E0000000020",
INIT_14 => X"0840024D810283021280400720C0348002854C001CC3158026A2040028090441",
INIT_15 => X"80901A0901A09018090188901A248054480C0C0041116DD0115E011599641E59",
INIT_16 => X"C6C8408514028028D06C0C5D20030BA1010021B000020402400501A090180901",
INIT_17 => X"4290C4290843908439084390843908439084390C4290C4290C4290C4290C4690",
INIT_18 => X"290C4210E4290C4310A439084310A439084310A4390C4290C4290C4290C4290C",
INIT_19 => X"5D54AAB556AA9556AAC310A439084310A439084310A439084210E4290C4210E4",
INIT_1A => X"0820825103A1600054C0F4012492490300C78C706428A1411133586294020A90",
INIT_1B => X"D4EA753A9D4EA753A92492492492492492492492492492492492492482082082",
INIT_1C => X"8086A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A353A9",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE024",
INIT_1E => X"5421EFAAFFD54AAF7D168B45AAAABDF5500002AA100000000000000000000000",
INIT_1F => X"043DF45FFD168AAA0855420AAAA843DFFFAAD1554005D7FD74AAA28400155005",
INIT_20 => X"2AA955FF5D003FE10F7803FEBAFFD5420AA080400155AAD5554AAF7802AB4500",
INIT_21 => X"AA8028B45A2AE82155A2FBFFEBA0800021550855555FFAA84001FFAAAE80010A",
INIT_22 => X"0085168ABAFFFBD54BAAAAE97400A2FBC20AAA284175EF55517DF555D2EBFE00",
INIT_23 => X"55AAAA954AA5D7FFFF45AAAA975EF007BD7555FFFBFDF55AAFBD55EF5D2EBFE1",
INIT_24 => X"BEFAAD1575EFAAAE974AA5D00175555D0015410F7AAAAAAA55043DE00FFFFD55",
INIT_25 => X"00000000000000000000000000000000000000000004174105D517DF55AAAAAA",
INIT_26 => X"D54AABC04001C51551471D7AAF1D05D2EBD56DB7DBEAEBFF551C042AA101D000",
INIT_27 => X"B50492EB842FB5508043FF55EBD56ABD75D5B470AABE8A3AFD7A2DF55400557F",
INIT_28 => X"8E82557FD2082000BEAE905C755003FE28E3D17DEAAEBDF40002550F47155AAD",
INIT_29 => X"5517DF40552ABDF45B6AEAFFD5F7A48017DAAFFFAE821C0A0717D1C5B575FFB6",
INIT_2A => X"F7D5C55D7492E90E3808756DA92EBFFD74BAE3AE85480FFFFC00AABE8E105C75",
INIT_2B => X"241043AE10EAF5C5547FF80954AA5D7FFAF7DA2AE905EF0075D5545E3F5EFF57",
INIT_2C => X"105D5B7FF7DB6AAAABC7BEDB505EFBEF5C7092FF801756D490A10438EBA4B8E9",
INIT_2D => X"F555D0028A00510000000000000000000000000000000000000000000000E124",
INIT_2E => X"8B45AAFBD54005D7BD54AAF78002155515157555AAD142040A2D57FFFFFFAEBF",
INIT_2F => X"DC01051AE955F7AAFBC0000AF843FF5500003FF55AAFD6AB455157D74BAF7AAA",
INIT_30 => X"E955FF557BD74EFFBACD41577B8400010F7AA8215555003FEAAAAC53DEB8A2FD",
INIT_31 => X"FEC20BAF7AA8015558517FF555D2ABDF51F782BCB47ABAE801FFAAFBEAA105D2",
INIT_32 => X"8554214FA2D3EAF57AFFDD7555082AA0AAA00557FEA8A2FDD64BAAF8282012AF",
INIT_33 => X"082A820AAAB842AA00000028AB0AAFF48547AE04174BA557BEABEFA2AA951FF8",
INIT_34 => X"0000000000002A80010557BFDFFFF7822A955FFFFC21FFF3BE40412DE02955FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000800000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303000048B3532C82D04A16002",
INIT_01 => X"210399800808004C1C20650E1E104368403008418984014902030006A8910200",
INIT_02 => X"480108A200000000444148E41E80F00A4104311868200200080000000988A390",
INIT_03 => X"0CA08220080000D004260A0240109028270012603000000030808C4208C000F0",
INIT_04 => X"4403A609A055306BC2C0735810CEE5100A0A48E16B8370E3808241D03845D002",
INIT_05 => X"ECE8698800791403AD3038AE079059A790E245A19A41E4120BAB86C00001D312",
INIT_06 => X"23208806000C3D220023C0021A21008891048C00040341121661E3C10000A064",
INIT_07 => X"0008045000220440000000090800102118400204A04100F040018019004B8001",
INIT_08 => X"0E11400810906441123323C0424190880B0108002000000880810F9002041200",
INIT_09 => X"22003C2309671584786E0F5A88889031EF9F05D884794FA03A24781810106D02",
INIT_0A => X"0409400E4282A00142400004DC3C82400702003200872003FB14080828400010",
INIT_0B => X"F050C3C00095000C008135040002010100800040001400C00401208800F01A14",
INIT_0C => X"08000002E0100000000800000220100000000800000001C87261C51C42390240",
INIT_0D => X"0400000280100000000800000360100000000800000035100040000000000000",
INIT_0E => X"00000000000004000000D8008000000000000001000000155000080000000000",
INIT_0F => X"000040000120EC00004002214000008000000000000200000000000094100040",
INIT_10 => X"001000000200050C000200000000000040080005800008000001000168000040",
INIT_11 => X"000800000000004008000448000040000000000001003C000008000008000D00",
INIT_12 => X"800800000000800000000001000008000017000100000000000010200002C800",
INIT_13 => X"150F5E0400101000227200800E271E00288400800208004C04C0080000000052",
INIT_14 => X"818082450000920280C544310041B408880EC51060461589225100063E9012D6",
INIT_15 => X"1410C3410C1410C1410C3410C100869A08618C00772201D899BA003591510A59",
INIT_16 => X"44E0110004480020986D4815044369A00006203041C3443043010C5410C3410C",
INIT_17 => X"0080001002008040100200800000060180000006008000100600804000020180",
INIT_18 => X"0000010060080201800000040100201802008040100201804000020180001006",
INIT_19 => X"64B261934D964C32698080401000000060080601800000040000201806008000",
INIT_1A => X"1451457A604C8D0C28A280CD145144C1863807E0500014385DAF345041488280",
INIT_1B => X"1A8D46A351A8D46A355555555555555555555555555555555555555545145145",
INIT_1C => X"1F60D068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D06A35",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE077",
INIT_1E => X"02ABFF087FFDF5508003FEBA087FD54BAAA84154005500000000000000000000",
INIT_1F => X"2EBFF5500003DF455555421EFAAFFD54AAF7D168B45AAAABDF55A2802AA10000",
INIT_20 => X"A843DFFFAAD1554005D7FD74AAAA840015500002AABA082E954005500021FF5D",
INIT_21 => X"FFD168BEF080028BFF0855555455500174BAA2AABDE0055517FF555555420AAA",
INIT_22 => X"0085168ABA0055574BA5555554BA5D0400155AAD1554AAF7802AB4500043DF45",
INIT_23 => X"AA5D0400010A2AA955FF55003FE10F7803FEBAFFD5420BA085168A00007BFDE1",
INIT_24 => X"1550855555FFAA84001FFAAFBEAB45002A97545F7D1555EF55043DF5555517DE",
INIT_25 => X"0000000000000000000000000000000000000000002A82155A2FBFFEBA080002",
INIT_26 => X"BFF55BC042AA101D0A28BC7007FFDF45080A3AEAA007BD2482BE84124285C000",
INIT_27 => X"4974004100021FF492AB8F7D1C0438E381451471D7AAFBD0492EBD56DB7DBEAE",
INIT_28 => X"557AFED1C5F470AABE8A3AFD7A2DF55400557FD54AABE84001C5550A28ABA142",
INIT_29 => X"B842FB5508043FF55EBD56ABD75D0428BEF005557545490012482B6A0BAE2849",
INIT_2A => X"557F6DA101475FDE10145F68A921C55504924955524AA140E0717DAADB50492E",
INIT_2B => X"F5D043AF6D405F78E3A1C2002000BEAA905C755003FE28E3803DEAAEBDF40002",
INIT_2C => X"7DAAFFFAE821C0A0717D1C5B575FFB6DF425575D7BEFB55002097555FFD5401E",
INIT_2D => X"010F784000AA5900000000000000000000000000000000000000000000020801",
INIT_2E => X"2000A2D57FFFFF7AEBFF55FF8028A00512EAAB45007FFFF55082EA8AAA087FC2",
INIT_2F => X"02155512AAAA085D04174100800021FF002EA8BEF5D0428ABA595557555AAFBC",
INIT_30 => X"402000FF802ABAA04552ABFF597FD74BAF7AAA8B45AAFBD54005D7BD54AAF780",
INIT_31 => X"2F955FFAAFBC0000AF843FF5500003FF55AAFD6AB4551002ABEF005555555000",
INIT_32 => X"A843DEB0A2FD5600051537DE005D557DE005D7BE8AA85555400100879560AA59",
INIT_33 => X"000417545FFD5421FF5D0428BEF0079FCABA598400010F7AA8215555003FEAAA",
INIT_34 => X"00000000000004001FFAAFBEAA105D2E955FF557BD75EFFBBCD415521FBFDF45",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000001000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB0A0791B1B41694368283C81F9996A091A32152007AB37B20E07C0C1E002",
INIT_01 => X"881FBC449030884C446A00000034824841280A00084000C8C212812EEA953231",
INIT_02 => X"C809AD5CB118E640A4F408FC011FF0002080000082CCC66609DB7DDDCB1F2036",
INIT_03 => X"4A100E4D3E4C90D290831C824A4204720B20048A88800000B8E0F91028C5500E",
INIT_04 => X"00144884922644001914830051110A71E03040F0105B001C662AE22DC08A3408",
INIT_05 => X"120340220B88820041CDC451B860A6506BEBD08265AE105714505F0152122449",
INIT_06 => X"207F7890752C037372A1D72A398CD084C890EA2950A37E270660182C0D2C8080",
INIT_07 => X"9378355E64B66F96231CC81D2DAB468D38C601C5FFF54FF1C9A46490261C4B39",
INIT_08 => X"7F105CAD1089654115814FC60284A1A93B46F4621030C800001D7FA56891162E",
INIT_09 => X"E00A003C832D25328526C082DF9AB88C104024C09639441807B78661090C24A1",
INIT_0A => X"4FD32A2E2A9992944AF2D611C3FC01B2152109204C28B67061EC928920C569E7",
INIT_0B => X"F0313FE92C22F21CA0B363C0A242502028901408154218144D712664A5F15AC1",
INIT_0C => X"B2F0F1E01BE53FE1F000BE0FC41BE53FE1F000BE0FC80020130841840308653F",
INIT_0D => X"C3CB7F041BE1BFE1F000BE0FC41BE1BFE1F000BE0FCD806FFFAF0AE83080E2AE",
INIT_0E => X"1A7806013879BAA78FC103FF5F1F12F0380231F0BF9E3F02A7FFD63669C0E008",
INIT_0F => X"483136F200A822CBACAB9DDEB7F9BC291F30180309A0F83FE2B87C7D006FFF9F",
INIT_10 => X"D1C6184131B7980DFFFC03F00003F01FB931E9C1DBF8A30C2098DBE2FF7F2320",
INIT_11 => X"F060703080E29F1B71E9F6427EFE901C0E004C72BEC95FEF64E4090626DF15B7",
INIT_12 => X"EFAC6DFC8C0312A0024B83F07F3991E9F21DFFFA0A3C0202B8776AC7A7C9CBFF",
INIT_13 => X"88F4C1C64044A264601144C5F1787E1C812A510885C56620590350ACD3A7D5B7",
INIT_14 => X"9054204DF56A974F92C3E20F24301300082C38C4184F10281204888298284616",
INIT_15 => X"A238CE238C8238CE238CA238CC11C6411C670C10EB4124C2B3923BF5C9710C59",
INIT_16 => X"276A11A03444922898494C5504008401230E71B3100C1634E3138C8238CC238C",
INIT_17 => X"5094650142511405194450942511425114450944519425114250144519405194",
INIT_18 => X"0944509465114251146501465014051944509445094051942501465014051940",
INIT_19 => X"2124B2DA6924965B4D5094450940519425014650142511425014450944519405",
INIT_1A => X"7DF7DF6FEFFCFDFD796ED1DCF3CF3DF6CE7F7B9DB7FF3A7E1FBC6DB7E8418A88",
INIT_1B => X"EEF77BBDDEEF77BBDDF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF",
INIT_1C => X"024F77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDD",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE056",
INIT_1E => X"5574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF80000000000000000000",
INIT_1F => X"D16AABAF7AAA8BFFAA802ABFF087FFDF5508003FEBA087FD54BA080415400555",
INIT_20 => X"AFFD54AAF7D168B45AAAABDF55AA802AA1000003FEBA00002AABA5D2EBFEBAAA",
INIT_21 => X"00003DE005555575EFA2D142145A2FFE8B45FF80001555D2E955FFFFD5421EFA",
INIT_22 => X"F5D7FC00BA5D5568AAAF7AAAAAAAAA802AABA082E954005500021FF5D2EBFF55",
INIT_23 => X"BAFFD5420AAAA843DFFFAAD1554005D7FD74AAAA840014500517FFEF007BEABF",
INIT_24 => X"4BAA2AABDE0055517FF555504154BAA2FBEAA105D2E97410FFD16AAAA5D2ABDE",
INIT_25 => X"0000000000000000000000000000000000000000000028BFF085555545550017",
INIT_26 => X"D24821E84124285C51574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7800",
INIT_27 => X"428A925D2AB8EBABEDB6AA92F7AAA8BC7B68A28BC70075FDF45080A3AEAA007B",
INIT_28 => X"2A925FFFFD1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0A38EBA1C0",
INIT_29 => X"100021FF492AB8F7D1C0438E38145B575EFA2DB45145B6F5EFB6DF78E0514555",
INIT_2A => X"55517DFC70875EABC7557FC20AA415F68AAAF7AAAAA82BE8A28A921424974004",
INIT_2B => X"0FFDB6FABA542ABAE2AF7DF470AABE8A3AFD7A2DF55400557FD54AABE84001C5",
INIT_2C => X"EF005557545490012482B6A0BAE2849043AFED1C0E10492B6FFEFA105D2A9541",
INIT_2D => X"E005D2AAABEFFB8000000000000000000000000000000000000000000000428B",
INIT_2E => X"FF55082EA8AAA087FC20105504000AA5955554BAFFAEBDE10F7FBFDEBA007BFD",
INIT_2F => X"28A00512AA8AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3AAAAB4500557",
INIT_30 => X"57FFEFFFAA97545552A821EFFBD557555AAFBC2000A2D57FFFFF7AEBFF55FF80",
INIT_31 => X"AAAAA005D04174100800021FF002EA8BEF5D0428ABA597FD55FFA2FFD5555FFD",
INIT_32 => X"D7BD54AAF7800015551517DF45005168B55557FC0012087FEAABAF7AAAAA10F3",
INIT_33 => X"FFFFFFE005D2A95410F7FFFFEBA5D2EA8ABAFBFFD74BAF7AAA8B45AAFBD54005",
INIT_34 => X"000000000000002ABEF005555555000402000FF802AAAA04452ABFF592E80010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000006000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C030028180004003220200403302301C0381A0082",
INIT_01 => X"A74041C838394848188160000C42426041000000090800090210000008510200",
INIT_02 => X"080108200C1000004465580000C0080100000000010432400800800009882050",
INIT_03 => X"080200010C234040842248600210812183806584488000103080014E88C10000",
INIT_04 => X"0040584288A6C210003120000000001002A0E8A910A072101000400A00203040",
INIT_05 => X"04096A019400C118414A00014000002014100128005004020010A0C044C02800",
INIT_06 => X"20200A301223FC029931E9931900002224240249A6D3E808D51FE00909108222",
INIT_07 => X"0008040000220001820000010C0810211A440014A040200E8240089000080002",
INIT_08 => X"0040081A08944010007FA038020080880B0104182000000000090F8102041320",
INIT_09 => X"17E2FD200240B4A409223F020888100808200450001A401BF82C21185C81744A",
INIT_0A => X"0602A0244285180542402180D001BE1907939120000020044184890800011000",
INIT_0B => X"0F0400091081190E4490A502D2A36951B428DB14A688051A5E21214601A01A22",
INIT_0C => X"455D0018101480000000A01034101480000000A01033A0081300000000001880",
INIT_0D => X"0001A0F4101480000000A01034101480000000A0103142000040000000000000",
INIT_0E => X"00000000000041E8002900018040000000000000466800C20004090000000000",
INIT_0F => X"0000034D242C2000502000000080028000000000000000240946800142000040",
INIT_10 => X"20900000001A60F0000200000000002007F000322010480000000D1A00040440",
INIT_11 => X"2018000000000025D00008958010440000000000403F4000808800000068D240",
INIT_12 => X"101280008200800000000000086670000CC0000100000000000087C000301400",
INIT_13 => X"C8B5800720849A72700094A2202301F05103202420000810C219500150002800",
INIT_14 => X"81088A454110030212C140813204D0A0888C000118471DE126805432A62A1586",
INIT_15 => X"4096C4096C2096C2096C6096C444B6004B600C446B0104D09190013589701C11",
INIT_16 => X"108D19D1804A8000904C421852240821978221B0044245B25B456C0096C0096C",
INIT_17 => X"69DA368DA1695A568DA3685A1695A768DA3685A569DA768DA1685A569DA76C5A",
INIT_18 => X"85A569DA1685A369DA5695A368DA169DA7695A168DA3695A5695A368DA3695A5",
INIT_19 => X"7638C31C71C718638E685A569DA7685A368DA5695A768DA1685A7695A168DA36",
INIT_1A => X"1C71C73B676CEDED7DE2F4DDF7DF7DF7CE7F8FF0F4FA957FCF9F7CF7F40A0010",
INIT_1B => X"FE7F3F9FCFE7F3F9FC71C71C71C71C71C71C71C71C71C71C71C71C71C71C71C7",
INIT_1C => X"2BE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"0000000000000000000000000607C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF019",
INIT_1E => X"43DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFF80000000000000000000",
INIT_1F => X"D17DEBA0855421455555574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF8",
INIT_20 => X"87FFDF5508003FEBA087FD54BA000415400550428AAAAA84021FF007BD54BAAA",
INIT_21 => X"F7AAA8BFFAAD1554BA002A95555A28417400AAFBE8ABAF7FFD54AAAA802ABFF0",
INIT_22 => X"0FFFBD5545080417555A2D17FE1000003FEBA00002AABA5D2EBFEBAAAD16AABA",
INIT_23 => X"FFFFD5421EFAAFFD54AAF7D168B45AAAABDF55AA802AA100000001EF087FEAA0",
INIT_24 => X"B45FF80001555D2E955FFFF843DEAAA2803DFEF0855401FF082EA8B555D7FC21",
INIT_25 => X"00000000000000000000000000000000000000000055575EFA2D142145A2FFE8",
INIT_26 => X"6FA92552AB8FEFF78E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FF800",
INIT_27 => X"E001EF147BD2482BED57AE921451421555551574BAB68A2DA00FFFFFFE38085F",
INIT_28 => X"FFD24BAB68A28BC70075FDF45080A3AEAA007BD24821C04124281C0E2DA82BE8",
INIT_29 => X"D2AB8EBABEDB6AA92F7AAA8BC7B6D5524AA14209557DA28E15400BEF1EFA92FF",
INIT_2A => X"5D0E071FF0071EDA38F7F1D5555000417545B6D178E281C0A38EBA1C0428A925",
INIT_2B => X"70824A8B555C7FC2147F7D1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA10",
INIT_2C => X"EFA2DB45145B6F5EFB6DF78E05145552A925FFFF8E3DE82BE8E38FFF0851401C",
INIT_2D => X"000557FE8A00F38000000000000000000000000000000000000000000005B575",
INIT_2E => X"DE10F7FBFDEBA007BFDE005D2AAABEFFBAABDFEFAAFBC00BA007BC0000FFD542",
INIT_2F => X"000AA592ABFE00F7AA821FF557FC0010F7D168A105D55421455155554BAFFAEB",
INIT_30 => X"E95410F7D57DE00FFFBC00AAFBAAAAB4500557FF55082EA8AAA087FC20105504",
INIT_31 => X"2AA8AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3D5400BA5504155EFAAA",
INIT_32 => X"7AEBFF55FF8028A00512E975FF08557FEAAF7D157545080417545F7D56AAAA59",
INIT_33 => X"F7AAAABEF005542155000028B555D7FC2145F3D557555AAFBC2000A2D57FFFFF",
INIT_34 => X"0000000000007FD55FFA2FFD5555FFD57FFEFFFAA97545552A821EFFBAABDE00",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000004800000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992006",
INIT_01 => X"A34009C0383848481C00E0000E01426040000000080000080200010000510204",
INIT_02 => X"4801082048100000446558000080000041000000000622400800000009000010",
INIT_03 => X"080001038CA14840842248400210812102000400088000003080014688800000",
INIT_04 => X"000040048106000040120000000000100220C8A5108032140004500800603000",
INIT_05 => X"04096A009000410041480081000000201000012800400022801080C0C0C82000",
INIT_06 => X"232086381A8001220021E0021803002224240248040360889100100909000222",
INIT_07 => X"0008055000220409020000090C0810211A04001420602000D2500810000C4903",
INIT_08 => X"8040491A809041100001400042409098090006102000000000010F8102041320",
INIT_09 => X"340C013102002420012200820D89140800004010900A4010002C8118D0024412",
INIT_0A => X"A221A5000800914000400888C00100200B0310200008B2066313894800631400",
INIT_0B => X"0010000800010004088105020100008000400120800000200404002450004000",
INIT_0C => X"4409081C1000000000F001F02C1000000000F001F021141A12000000000010B0",
INIT_0D => X"383480CC1000000000F001F02C1000000000F001F023420000000004C3201C51",
INIT_0E => X"00019860078641084039000000000002C0E00E0E404900E200000000000B0380",
INIT_0F => X"120C8908146000105120000000000004004160C0301D07001D04820342000000",
INIT_10 => X"000021908C4842FC000000030F000FE00600103BA0000010C8462414E8000006",
INIT_11 => X"000004C3201C60A400100DD5800000013098038D40309D000000C2419120A740",
INIT_12 => X"901A800030040902C0807C0E00C440100DDD000000411C81078884004035DC00",
INIT_13 => X"140A000410401400201020820022000250400040002211148019064200402A32",
INIT_14 => X"01889A4543148282A01415B04009904A80890033679459A926801054001C0050",
INIT_15 => X"159201592055920559205592070C901AC901A100804000801210541403C05130",
INIT_16 => X"2460010004428008904C085D44200D8001112804CDE1C483480D201592015920",
INIT_17 => X"0080200806008020000000004000020080200802000000000000000008020480",
INIT_18 => X"1000008020080000000000020080200000000000080600802008000000400000",
INIT_19 => X"5841040002082080000180200000000020180200800000000100200802000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000005428A94",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"E480000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE031",
INIT_1E => X"BC00AAF7D5575455D557DFEF002AAAB55002E820AAAA80000000000000000000",
INIT_1F => X"AEAAB55007FD74AAAA843DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFF",
INIT_20 => X"2802AA10FFFFFDE0008556AABA5D2ABFFEFFFAAAAAAAF7D57FFEFF7D555555A2",
INIT_21 => X"085542145552ABDFEFFFAA801EFFFFBFDF550000175555504175450055574AAA",
INIT_22 => X"0082A975EF00003DF55555168A00000428AAAAA84021FF007BD54BAAAD17DEBA",
INIT_23 => X"AAFF802ABFF087FFDF5508003FEBA087FD54BA000415400557BD74BAFFD14000",
INIT_24 => X"400AAFBE8ABAF7FFD54AAAAAEA8ABA55557FEAAA2843FF55A2AEA8B55AAAABDE",
INIT_25 => X"00000000000000000000000000000000000000000051554BA002A95555A28417",
INIT_26 => X"C20825D7FE8A92FFFFC70BAE3D155555415178FD7082EAAB550820870BAAA800",
INIT_27 => X"578FFFEBD55557DBEA4AFB550871D7482AA8E3DFFFAAFFD04AA415B52492B6F5",
INIT_28 => X"0E175550051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7A0ADABAEBD",
INIT_29 => X"47BD2482BED57AE921451421555524BDFD7FFA4801D7F7F5FDF55000E1754541",
INIT_2A => X"1C7BD2482E3D1450381C20905EF08003AF55415F6DA38080E2DA82BE8E001EF1",
INIT_2B => X"5BEAAAFB55ABA0BDE02EB8A28BC70075FDF45080A3AEAA007BD24821C0412428",
INIT_2C => X"AA14209557DA28E15400BEF1EFA92FFFFD24BAB6A4A8A82495F78E92AA843DF4",
INIT_2D => X"B450800174BAA680000000000000000000000000000000000000000000055524",
INIT_2E => X"00BA007BC0000FFD542000557FE8A00F3FFD54BAAAD15754508556AB45002AA8",
INIT_2F => X"AABEFFB803DEAAAAD56ABEFAAD5575EFF7803DF45085557410AEAABDFEFAAFBC",
INIT_30 => X"57FF55082E97555002E955550C55554BAFFAEBDE10F7FBFDEBA007BFDE005D2A",
INIT_31 => X"2ABFE00F7AA821FF557FC0010F7D168A105D554214551003FF45FF8400145FFD",
INIT_32 => X"87FC20105504000AA597FC2010A2D1554AA5500021EF000028B55087BFDEBA04",
INIT_33 => X"007FE8A00A2803FF45F7AABDF55AA843FE10AEAAAAB4500557FF55082EA8AAA0",
INIT_34 => X"00000000000055400BA5504155EFAAAE95410F7D57DE00FFFBC00AAFB8028A00",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"A140084000080048040100000202026040000000180800080200010048510204",
INIT_02 => X"080108000090000004655C000080000051000000000402400800000009000010",
INIT_03 => X"0000000100300C40842240000210810002800584488000103080894288800000",
INIT_04 => X"0002584280A2C21000110300100000100220C8C910A032541000090A00643000",
INIT_05 => X"04092A001400D100410A002140004020140001A9005000004810A1C0044D2800",
INIT_06 => X"0360000010EFFD229911C9911820002080258A09A2D3E102137FE0094910A222",
INIT_07 => X"0000004000220400120000090C0810210A040034A040000046180810000C4907",
INIT_08 => X"80404050D88C24510001400042008088090004012000000000010F8102041320",
INIT_09 => X"20080120024030A4090200828C880208002044C0843B44100228A1585C81740A",
INIT_0A => X"142180860A84802042C82180D0010039039390200008B20E2300086800400640",
INIT_0B => X"003000091084190644810502D0A16850B4285B14A688011A1409212008F05E20",
INIT_0C => X"400104080010001E0FF00010000010001E0FF0001002200A1300000000000080",
INIT_0D => X"000080000010001E0FF00010000010001E0FF000100440000040F517CF600000",
INIT_0E => X"E587F9E000004008100800008000ED0FC7E000004000804000000809963F1F80",
INIT_0F => X"36000100202C0020100000000802419660CFE7C0F00000000800810040000040",
INIT_10 => X"0618E7B0000800000003F80FFF0000200018021000030C73D80004000000585F",
INIT_11 => X"078A8FCF600000201802008001006AA3F1F80000400000000B0BD6C000200000",
INIT_12 => X"0041120370DCAD1FC18000000040180200800005D5C3FD800000806008100000",
INIT_13 => X"48A480072284983230101402200200111103202420000880C218000150100800",
INIT_14 => X"2B888A4500048240C08400843204502000890001000415E12480003002944281",
INIT_15 => X"0480004800048000480004800004002240020854884000901212140011C01079",
INIT_16 => X"346D19D1A4C08028904C4E1D7224086590800420044040020004004480004800",
INIT_17 => X"68DA368DA368DA368DA368DA368DA1685A1685A1685A1685A1685A168DA36CDA",
INIT_18 => X"8DA3685A1685A1685A1685A368DA368DA368DA3685A1685A1685A1685A1685A1",
INIT_19 => X"40000000000000000068DA368DA368DA1685A1685A1685A1685A368DA368DA36",
INIT_1A => X"3CF3CF6FE23CCD8D00A281F5B2DB2CA78A543EBC57A10A245DA975D640088884",
INIT_1B => X"3E1F0F87C3E1F0F87CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"5DA9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0F87C",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00B",
INIT_1E => X"40000000043DF55087BC01EF007FD75FFFF84000AAFF80000000000000000000",
INIT_1F => X"2EBFE10A28028AAAAAFBC00AAF7D5575455D557DFEF002AAAB55002E820AAAA8",
INIT_20 => X"2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFAA95545552ABFE00087BC00AA08",
INIT_21 => X"007FD74AAAAD57FF45002A975FF007BE8BFFA2FBFFFFFAAD5400AAFF843DFEFA",
INIT_22 => X"5AAFBE8A00082A97410F7D5555EFAAAAAAAAAF7D57FFEFF7D555555A2AEAAB55",
INIT_23 => X"450055574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFFAA8200055555554",
INIT_24 => X"F55000017555550417545000015545087BC2010AAD54014500516ABFFA2AABDF",
INIT_25 => X"0000000000000000000000000000000000000000002ABDFEFFFAA801EFFFFBFD",
INIT_26 => X"AAB550820870BAAA8407000140038F450075C71FF087BD75D7FF84050BAEB800",
INIT_27 => X"AB8E10007FC50BA002ABFE00AA8A2AABABEFFC70BAE3D155555415178FD7082E",
INIT_28 => X"DB45082EB8E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFA497545552",
INIT_29 => X"BD55557DBEA4AFB550871D7482AAD17DF451C24955EF0875EFBD7B6F1FFFC7BE",
INIT_2A => X"F7AA87000415B5057DAAFBE8A10082092410EBD5505EFB6A0ADABAEBD578FFFE",
INIT_2B => X"D005B6ABC7B6AABFFED0051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEF",
INIT_2C => X"D7FFA4801D7F7F5FDF55000E17545410E17555000E17545007BC0000BED14217",
INIT_2D => X"555F784174AAA280000000000000000000000000000000000000000000024BDF",
INIT_2E => X"754508556AB45002AA8B450800174BAA684174105D042AB550055555FF007BD7",
INIT_2F => X"E8A00F384175555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7FFD54BAAAD15",
INIT_30 => X"57DF55FFD57DF55FFFBD5400A2AABDFEFAAFBC00BA007BC0000FFD542000557F",
INIT_31 => X"803DEAAAAD56ABEFAAD5575EFF7803DF45085557410AED17FF455D04155FF005",
INIT_32 => X"07BFDE005D2AAABEFFBAE97410087BC21EFA2FFEAA00000002010A2D5421FFFF",
INIT_33 => X"087BC0010FFD1401EF087FE8B55FFAEBDFEF0855554BAFFAEBDE10F7FBFDEBA0",
INIT_34 => X"000000000000003FF45FF8400145FFD57FF55082E97555002E955550C2E95555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000002000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000006",
INIT_01 => X"0000098218302849180060000C004260413C0A61590001D90213C80000110200",
INIT_02 => X"680108220010000054400C00008000004100000001200240080080000908A011",
INIT_03 => X"000A0000040020400002021000000008428065044880001030818C0008C10000",
INIT_04 => X"00005042882A8210003000000800001000806080100040140080040800003140",
INIT_05 => X"0400000840000098410800010001002000000000004000002010000040002000",
INIT_06 => X"03600810100001220911E0911902000020200200A253E8000C0010080800004C",
INIT_07 => X"000408C0002204400200000B080000010C040004A0400000C0000810000C5901",
INIT_08 => X"000008002A84300000014000C2008088090008002000000000030F8000001220",
INIT_09 => X"0008012100000200001200820888010800200000000840100028800004801440",
INIT_0A => X"000090220000040400480000D0010009049090200008B2022384800802010000",
INIT_0B => X"001000090001090A4C81240050A328519428CA14328C840A5820000101500400",
INIT_0C => X"00510008100400000000A00000100400000000A00000000A12000000000000B0",
INIT_0D => X"00012000100080000000A00000100080000000A0000540000000000000000000",
INIT_0E => X"00000000000000A8000900010000000000000000060000420004000000000000",
INIT_0F => X"0000024000240000102000000080000000000000000000240000800140000000",
INIT_10 => X"0080000000120CFC000000000000000001280013E010000000000900F8040000",
INIT_11 => X"2000000000000001480006D5801000000000000000091F0000800000004807C0",
INIT_12 => X"901A800080000000000000000820080006DD000000000000000002A00019DC00",
INIT_13 => X"0200800522C01252501086222082000010012024200000048019502000000C32",
INIT_14 => X"0080004501000200089400005200D0820008000000104C4800010600BC228404",
INIT_15 => X"0001040010000104001000010440080000822900000000801010500A13404111",
INIT_16 => X"32851951A0CA8080924C06403600086491900224002200400440104001040010",
INIT_17 => X"284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A128CA328CA",
INIT_18 => X"84A1284A1284A1284A1284A328CA328CA328CA328CA328CA328CA328CA328CA3",
INIT_19 => X"10000000000000000028CA328CA328CA328CA328CA328CA328CA1284A1284A12",
INIT_1A => X"69A69A250B61004055CD1439248209070CCCF48DE68A8900401038E2550A0010",
INIT_1B => X"341A0D068341A0D068A28A28A28A28A28A28A28A28A28A28A28A28A29A69A69A",
INIT_1C => X"56C1A0D269341A0D068349A4D068349A4D068341A0D269341A0D269341A0D068",
INIT_1D => X"0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE052",
INIT_1E => X"57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D00000000000000000000",
INIT_1F => X"D1575EF00557DF555D040000000043DF55087BC01EF007FD75FFFF84000AAFFD",
INIT_20 => X"7D5575455D557DFEF002AAAB55002E820AAAA843DFEF00517DEBA007BFDFEFFF",
INIT_21 => X"A28028AAAAAAABDF45F7803FFEF555568AAAF7802AA00FFFBD7555087BC00AAF",
INIT_22 => X"5087BD54BA550417400085155555082A95545552ABFE00087BC00AA082EBFE10",
INIT_23 => X"555D043DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00AA552E9554",
INIT_24 => X"BFFA2FBFFFFFAAD5400AAFF8402000A2FFFDF555D7BE8BFF5D51575EFA280175",
INIT_25 => X"000000000000000000000000000000000000000000557FF45002A975FF007BE8",
INIT_26 => X"D75D7FF84050BAEBDF78F45B68010482415B471C7E3DF451EFBEFBFAF4549000",
INIT_27 => X"17DE82007FFAFEFE3DB505EF1C5B7AF45490407000140038F450075C71FF087B",
INIT_28 => X"FFD55451C7FC70BAE3D155555415178FD7082EAAB550820870BAAA8438FFF005",
INIT_29 => X"07FC50BA002ABFE00AA8A2AABABEAEB8F45F78A3DFD741516DAAAE38E2DA28EB",
INIT_2A => X"FFFFC20BA5D2E905550071D54825D0A1543808515756D1C2497545552AB8E100",
INIT_2B => X"F5D55505FFBE801256D490E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92",
INIT_2C => X"451C24955EF0875EFBD7B6F1FFFC7BEDB45082EB8002000AAFFFDF6D417FEABE",
INIT_2D => X"5EFF7FBE8B5500000000000000000000000000000000000000000000000517DF",
INIT_2E => X"AB550055555FF007BD7555F784174AAA2FBEAB45F78402010007BD5545AAFFD5",
INIT_2F => X"174BAA68028BEF00517FE10007BE8BFFAAFFC01FF557FE8B550004174105D042",
INIT_30 => X"57FEAAAAAEBFEAAAAFFD5545557FD54BAAAD15754508556AB45002AA8B450800",
INIT_31 => X"04175555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7AAAAB45F7AEBFF45085",
INIT_32 => X"FD542000557FE8A00F3FFC00BA552E80145005557400552A954BA0051575EF55",
INIT_33 => X"A2FBFDFFF007FE8BFF5551401EFF784021FF002ABDFEFAAFBC00BA007BC0000F",
INIT_34 => X"000000000000517FF455D04155FF00557DF55FFD57DF55FFFBD5400A28400010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000004000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A14009801830084C182060000C10424840000000080000080200000000110204",
INIT_02 => X"0801080200100000046558040080000041000000002402400800000009008010",
INIT_03 => X"00020201040000D0842242024210810802006400088000003080054288C10000",
INIT_04 => X"0000400088020000003020002000001002A0E881108032100002000800203040",
INIT_05 => X"04092A081000411841480001000000201000012800400010001081C040402000",
INIT_06 => X"03600810100001220001E0001802002020240208000369001500100909000266",
INIT_07 => X"0000004000220440020000090C0810210A040004A0410000C0000810000C4901",
INIT_08 => X"0040480000802100100140004200808809000C002000000000010F8102041320",
INIT_09 => X"2008012000000000000200828888800808000410800840100220211850004442",
INIT_0A => X"040180240A80800442400004C0010000060210200008B2022304880800010000",
INIT_0B => X"0030000000010008008020020100008000400120800004004821202001A05A00",
INIT_0C => X"40510008101480000000A01004101480000000A0100000001300410402080080",
INIT_0D => X"0001A004101480000000A01004101480000000A0100540000040000000000000",
INIT_0E => X"00000000000040A8000900018040000000000000460800420004090000000000",
INIT_0F => X"0000034000082000102000000080028000000000000000240800800140000040",
INIT_10 => X"20900000001A00000002000000000020013000100010480000000D0000040440",
INIT_11 => X"2018000000000021500000800010440000000000400900008088000000680000",
INIT_12 => X"000000008200800000000000086010000080000100000000000082C000100000",
INIT_13 => X"000080000004924040008020000200101100004000000000C019500050000800",
INIT_14 => X"2B088A4541008240001000804000108280800001001051A12481041080801010",
INIT_15 => X"4480004800048004480044800044000240022100884000901210440003C14110",
INIT_16 => X"06E00000044200009849485D4020080000140004046240020044000480044800",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802000000400",
INIT_18 => X"0000000000000000000000020080200802008020080200802008020080200802",
INIT_19 => X"1000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"1451451AA654199951A24454514514F0CA940FE0D39712615FAD555204428290",
INIT_1B => X"CA6532994CA65329945145145145145145145145145145145145145145145145",
INIT_1C => X"670E572994CA6532994CAE572B95CA6532994CA6532B95CAE572994CA6532994",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE01C",
INIT_1E => X"03FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF0800000000000000000000",
INIT_1F => X"7FFDF45FFFBC2010AAD57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D0",
INIT_20 => X"0043DF55087BC01EF007FD75FFFF84000AAFF8002155AAFFE8B45AAD54000008",
INIT_21 => X"00557DF555D517FEBA082A801EFF7FBD5400FFD568B555D00155EF0804000000",
INIT_22 => X"AF7FBFDE00A2FBC0145005168A10AA843DFEF00517DEBA007BFDFEFFFD1575EF",
INIT_23 => X"EF5D7BC00AAF7D5575455D557DFEF002AAAB55002E820AAAA803FEBA082AAAAA",
INIT_24 => X"AAAF7802AA00FFFBD7555082E82155FFAEAAB55AAD568B455D00154BAFFFBD75",
INIT_25 => X"0000000000000000000000000000000000000000002ABDF45F7803FFEF555568",
INIT_26 => X"451EFBEFBFAF4549003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC700000",
INIT_27 => X"5EDB6DAADF470280075FFF45E3F1C7038A2DF78F45B68010482415B471C7E3DF",
INIT_28 => X"0A175C7000407000140038F450075C71FF087BD75D7FF84050BAEB8002155BEF",
INIT_29 => X"07FFAFEFE3DB505EF1C5B7AF45495B7DEAA0824851EFEBFBD2410EBD168B7D41",
INIT_2A => X"AA8038EAA0824A8AAAEBF5FAE28AAF1C2155005F68A10A28438FFF00517DE820",
INIT_2B => X"D4104104AAF7F1D75EF557FC70BAE3D155555415178FD7082EAAB550820870BA",
INIT_2C => X"45F78A3DFD741516DAAAE38E2DA28EBFFD55451C2087155EBA4A8B7DAADF68B7",
INIT_2D => X"FEFA2AEAAB55000000000000000000000000000000000000000000000002EB8F",
INIT_2E => X"2010007BD5545AAFFD55EFF7FBE8B5500043FE00F7D17FEBAA2D5574BAAAD17D",
INIT_2F => X"174AAA28002155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAB45F7840",
INIT_30 => X"BC2000AAD16ABFF002A975450004174105D042AB550055555FF007BD7555F784",
INIT_31 => X"8028BEF00517FE10007BE8BFFAAFFC01FF557FE8B55007FFDEAA0004175FFA2F",
INIT_32 => X"02AA8B450800174BAA68428AAA08042AABAAAD56AABAAAD140155087FEAA10A2",
INIT_33 => X"A2842ABEFAAFBE8BFF0004020AAFFD5555EF557FD54BAAAD15754508556AB450",
INIT_34 => X"0000000000002AAAB45F7AEBFF4508557FEAAAAAEBFEAAAAFFD5545550015555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000047FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B83008481800E0000C26426040000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"00080D4912E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"000048048002400048150000000002504230C899109032100020160880223000",
INIT_05 => X"040B2A229100410041088011100022201200012840440000B01088C0005C2400",
INIT_06 => X"03286A287E4003225021C5021880C02000A40249048363A5990010090908022A",
INIT_07 => X"8320694044222987020C80152D8910210A0400252B74200045C86810000C5B05",
INIT_08 => X"00404126509804400501400242C0B0B83B0134702000000000191FA162841324",
INIT_09 => X"2008013002000220001240820F8B2A08000040409018401001200159D80D64AA",
INIT_0A => X"91019B02080885200042E098C00101B0070310200008B60A23A51B2802067327",
INIT_0B => X"003000080802500C088325828102408120409120940680100504022148504440",
INIT_0C => X"1501D5761B011986695014A96E1A8119865A5018C5A0A00012004104020808B0",
INIT_0D => X"A2600AAE1A811986695014A96E1B0119865A5018C5AF0062C38A4DB680A0D824",
INIT_0E => X"1DB528802CAB184E8F4101621B1BAC845542056A289A1BB2078A922DA2A8B180",
INIT_0F => X"7A3D94392000224ACDE215883078681B5C05AA429189B60AC43CEC7F0272C384",
INIT_10 => X"134CD551BCA1C90006C0C2958502861120C003104289A668B8CAB27010633831",
INIT_11 => X"82806CA64090B89E015AAA880E48382EB8804B020A06020C67061BC785938085",
INIT_12 => X"470126C6284B2D20410AB4503089C00A8280819A5539D503336D61056ABA0062",
INIT_13 => X"000080060040142020015001004A00080042004000E8089C9003066E03513E41",
INIT_14 => X"010CBA45367082014000908020349320008000A1000C09A9348498B000000000",
INIT_15 => X"C32A0832A0C32A0C32A0832A0C19504195040040000000801010028001400010",
INIT_16 => X"2468118104400000904C0C0964200841010954000444D280140050C32A0832A0",
INIT_17 => X"4090240902409024090240902409024090240902409024090240902409024090",
INIT_18 => X"0100401004010040100401024090240902409024090240902409024090240902",
INIT_19 => X"0000000000000000004010040100401004010040100401004010040100401004",
INIT_1A => X"410410502A441495418984700000005088804180C0B10A04D0A7104201400284",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000010410410",
INIT_1C => X"7800000000000000201000000000000000000008040000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE060",
INIT_1E => X"4155EFAA842ABEFA280155EFFFFBC01EF0855400005500000000000000000000",
INIT_1F => X"FBFFF4508514000000003FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF080",
INIT_20 => X"280154BA5555401EFFFD5421EFA2FFFFF555D51575FFA2FFD75FF550015400FF",
INIT_21 => X"FFFBC2010AAD568AAAAAD142145FF80155EF0051555FF0804155FFF7D57DF45A",
INIT_22 => X"008001540008514215555003DFFFA28002155AAFFE8B45AAD540000087FFDF45",
INIT_23 => X"0000040000000043DF55087BC01EF007FD75FFFF84000AAFF802ABFFA2AABFE1",
INIT_24 => X"400FFD568B555D00155EF085168B45085142010FFAE800AA5D7BFDF45F7FFEAA",
INIT_25 => X"000000000000000000000000000000000000000000517FEBA082A801EFF7FBD5",
INIT_26 => X"7DF7DA2AEB8FC70000175EFB6802DBC7BE8A155EFE3FBC71FF145B4203855000",
INIT_27 => X"5D05EF550E15400E3F1FFF7D085B420381C003DE10BEF5EDAAAAAD547038EBD5",
INIT_28 => X"04105C7F7DF78F45B68010482415B471C7E3DF451EFBEFBFAF45495F575FFBEF",
INIT_29 => X"ADF470280075FFF45E3F1C7038A2DB68ABAB6D145145FF84155D7085B555C714",
INIT_2A => X"EB8428BEFBEA4BDE28140A1543800514515549003FFC7BE8002155BEF5EDB6DA",
INIT_2B => X"2417FFFF7DE3F1EFA10140407000140038F450075C71FF087BD75D7FF84050BA",
INIT_2C => X"AA0824851EFEBFBD2410EBD168B7D410A175C7005B6DB55145140000FFAE8508",
INIT_2D => X"5EF557BC20AA5D0000000000000000000000000000000000000000000005B7DE",
INIT_2E => X"FEBAA2D5574BAAAD17DFEFA2AEAAB550004175FFF7803DF45FFAE955EFAAFBD5",
INIT_2F => X"E8B55007FD75FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D043FE00F7D17",
INIT_30 => X"015555007FD5545550400145FFFBEAB45F78402010007BD5545AAFFD55EFF7FB",
INIT_31 => X"8002155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAAAAFFD555545FF8",
INIT_32 => X"07BD7555F784174AAA2842ABEFFF803DEAA5D2E974AA00515754500003FF55FF",
INIT_33 => X"555540000FFAE97410007BFFFFFA2D57FE105D04174105D042AB550055555FF0",
INIT_34 => X"0000000000007FFDEAA0004175FFA2FBC2000AAD16ABFF002A97545007FFFF45",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000004000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C048000C048400380000007024040000000080000088200002802153231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"421A0A0012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"02004000890200001837800001998C31C090609C104000102002140900003548",
INIT_05 => X"0402002BC200009841090001200006200800000020480010A4100100001C2000",
INIT_06 => X"033432287FC003230001D0001806C0060CB0622000037085C800100C0C200008",
INIT_07 => X"135038CE64B663DFA314C803292140890C0601F472D1640051F80C10020C493F",
INIT_08 => X"00000167C081000011814004C20481A92940EA7A3020480000071F846890162E",
INIT_09 => X"D40C01240008000080024082488BAF08000020000208401004300421800F04F8",
INIT_0A => X"F9F80FA0200E0BF40063FF9DC0010000180018200408B27E234913E900067F04",
INIT_0B => X"001100002002801000A04200000000000000000000029D204B7C0382FD0100F3",
INIT_0C => X"9628F97E0B348EDAC3900F6EFA0B158EDA93900F6EE230381208008001007A80",
INIT_0D => X"EAE64BCA0B158EDAC3900F6EFA0B348EDA93900F6EE8421392C96B1237E0D8BD",
INIT_0E => X"4CAEAD412EDD2B47CFF812A383430C669E622DBC31D73F6006A5891533EF9500",
INIT_0F => X"2E19B8BA30E022DAD8C100CA39E8CEBE66C2B083798D341B10DE7E14400392C7",
INIT_10 => X"32966471A9C5DD00B12728D5360234D62A49FAB442994B3238D4E2FB10463665",
INIT_11 => X"F0FABAC800DA550C29F36A8A2554E48A6430469392526208C6CC95C33717D885",
INIT_12 => X"2B416A51B60585A5C28895962502E9F36A828C4999AF580395542D27CDBA0020",
INIT_13 => X"0000800000001E404011F066000A000EE040000000873FB80B8A00EF03F56CC1",
INIT_14 => X"2284304D667C06CC6816B300403C13E2000000460010400000010CE080801010",
INIT_15 => X"872F0872F0C72F0872F0872F0C597863978421000800209010104ACA03414110",
INIT_16 => X"01000000104280009048004000000800001D5E05182493C5BC5AF0872F0C72F0",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0802008020080200802008000000000000000000000000000000000000000000",
INIT_19 => X"1000000000000000000080200802008020080200802008020080200802008020",
INIT_1A => X"492492240F010000146E502D4514510246088881360A95118B120CB054420210",
INIT_1B => X"6432190C86432190C82082082082082082082082082082082082082092492492",
INIT_1C => X"7FEB2592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2590C8",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"5421FF00042ABEFFF8400010082EAABFF55002ABEF0800000000000000000000",
INIT_1F => X"002ABEFFFFBD54000004155EFAA842ABEFA280155EFFFFBC01EF085540000555",
INIT_20 => X"AFBE8AAAA2D540000F7D57DF55A2AABFFEF08556AA10000028AAAFFD15541000",
INIT_21 => X"085140000005168AAA087BFFFFF5D04001FF00041554555557FE005D003FE10A",
INIT_22 => X"F0851555FF082AA8B55F7AEA8BEF5551575FFA2FFD75FF550015400FFFBFFF45",
INIT_23 => X"10AAD57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D0000145082E955F",
INIT_24 => X"5EF0051555FF0804155FFF7842AA100000020BAAA801541055042ABEFFFFBD54",
INIT_25 => X"0000000000000000000000000000000000000000005568AAAAAD142145FF8015",
INIT_26 => X"C71FF145B42038555F401D71C0A2DBC7EB80000280824ADBD7490E28BEF08000",
INIT_27 => X"A2DA82FFDB5243800002FBD7EBFBD24101C00175EFB6802DBC7BE8A155EFE3FB",
INIT_28 => X"5B7AE1041003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7005F6AA381C0",
INIT_29 => X"50E15400E3F1FFF7D085B420381C5B6AA82147FF8FEF410E001FF000E1755555",
INIT_2A => X"49000017D142E905EF1451525C7082AADB45F7AEA8BEF555F575FFBEF5D05EF5",
INIT_2B => X"041002FBEFEBFBD2410AADF78F45B68010482415B471C7E3DF451EFBEFBFAF45",
INIT_2C => X"BAB6D145145FF84155D7085B555C71404105C7F7842FA381C0A00082AA8A1041",
INIT_2D => X"F55002AA8BEF000000000000000000000000000000000000000000000005B68A",
INIT_2E => X"DF45FFAE955EFAAFBD55EF557BC20AA5D7BC01555D2EBFF55A284000AA08003F",
INIT_2F => X"AAB55007BE8AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D04175FFF7803",
INIT_30 => X"E821FF082A97555557FE8A0000043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AE",
INIT_31 => X"7FD75FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D7BE8A005D7FEABFF002",
INIT_32 => X"AFFD55EFF7FBE8B550004001FF5D2A801EF5D5142145082EBFF55F7AAAABEF5D",
INIT_33 => X"552A82010A2AA8000008043FFFFA2FBC2010A2FBEAB45F78402010007BD5545A",
INIT_34 => X"0000000000007BEAAAAFFD555545FF8015555007FD5545550400145FF843DEAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400986B830E84D182260000C1042684001000008220008A20019080A510200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00020201926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"00104884880A4400403003005800027102A0E8C110D83210642EA809C0203040",
INIT_05 => X"04092A08138041184109C001380000201A008128044E00754010C9C192D82400",
INIT_06 => X"032C7E201800012372A1D72A180000204024024954A3670819001009092C0222",
INIT_07 => X"0164004000220B40020C80052C0A12292A040005715540015E006810001C4B01",
INIT_08 => X"0040549032881001140140024200808839005C002010800000155F8122851320",
INIT_09 => X"6008012C80481284881280825A988008000040808629441005B3071859006442",
INIT_0A => X"0001B0200810940400720005C0030192072310200028B6022346080802E001A5",
INIT_0B => X"003000206822F20CA8826AC2A14250A128509528954404144C20042501004000",
INIT_0C => X"03D404A41AA5B7344C10B383081BA4B7341C10B3831034081200000000000430",
INIT_0D => X"5A2B2C381BA4B7344C10B383081AA5B7341C10B383110218CB0E54C2EA404A4F",
INIT_0E => X"3548B3A008E730A01AB113A5524E6ACA678001CE3E20A5B284ED1132909C7288",
INIT_0F => X"0A3C066430202021252991C22C99731014AC3CC0C0B8182597A801610218CB0C",
INIT_10 => X"A5C8825194332B018A444AEA2701288A15A151EC5952E44128CA194517354C18",
INIT_11 => X"635232D50048A411C158BB0A7910142C771804C8A0ADA2E6A983014780CA28B2",
INIT_12 => X"6E4023F8BE8E3E1E0109472C3EB50158BB02D09852745F80112C428562EE0353",
INIT_13 => X"00008002414032646000826080C20001104240480068001C9B9150A000029704",
INIT_14 => X"1118BA4510008241C80290882400908000A000A1000809A93485D61000000000",
INIT_15 => X"40000000000000040000000000000020000000040000008010122A8201410058",
INIT_16 => X"246A10A1044101A89A4D0C096420184321040002844840000000004000000000",
INIT_17 => X"5094250942509425094250942509425094250942509425094250942509425094",
INIT_18 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_19 => X"0000000000000000005094250942509425094250942509425094250942509425",
INIT_1A => X"75D75D7FEDFDFDFDFBEEF9DD555555F7EEFF3F7DF7FF3E7E1FBF7DF7E24502A8",
INIT_1B => X"FAFD7EBF5FAFD7EBF5D75D75D75D75D75D75D75D75D75D75D75D75D75D75D75D",
INIT_1C => X"7FEFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F780000000000000000000",
INIT_1F => X"AA97400AAD540155A2D5421FF00042ABEFFF8400010082EAABFF55002ABEF085",
INIT_20 => X"A842ABEFA280155EFFFFBC01EF08554000055043DEBAF7843FFFFF7AABDF55A2",
INIT_21 => X"FFFBD5400005568A1055043DEBAAAFFE8B45557FD7410552EAAABAAA84155EFA",
INIT_22 => X"AA2FFE8ABAAA8428A00087BD7555FFD56AA10000028AAAFFD15541000002ABEF",
INIT_23 => X"55A2803FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF085557545FFD17DEB",
INIT_24 => X"1FF00041554555557FE005D0000155557BEAABA5D2ABDF450851420AA5D7FD55",
INIT_25 => X"0000000000000000000000000000000000000000005168AAA087BFFFFF5D0400",
INIT_26 => X"ADBD7490E28BEF08516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EB800",
INIT_27 => X"03FFD7EBA4BDF45AAAA90410BEDF45155A2DF401D71C0A2DBC7EB80000280824",
INIT_28 => X"2AAFA82B680175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550E38E92EB8",
INIT_29 => X"FDB5243800002FBD7EBFBD24101C556FA38490A3FE92BEFFEAB45417FD24385D",
INIT_2A => X"00515056DE3D17FE92BEF1EFA92AA8428A10007FD557DFFDF6AA381C0A2DA82F",
INIT_2B => X"5085B400925D7FD557DA2803DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7",
INIT_2C => X"82147FF8FEF410E001FF000E17555555B7AE10410E00155497FEFABA4120B8F5",
INIT_2D => X"ABAA2FBD7545AA8000000000000000000000000000000000000000000005B6AA",
INIT_2E => X"FF55A284000AA08003FF55002AA8BEF00517FE00082EBDF45AA8428A10085568",
INIT_2F => X"C20AA5D2EA8A00A2803DF45AA843DF55AAAE82000F7FBD5545AAFBC01555D2EB",
INIT_30 => X"FE8B55087FC00BA552ABFE10F784175FFF7803DF45FFAE955EFAAFBD55EF557B",
INIT_31 => X"FBE8AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D517FEAA082EBFE10F7F",
INIT_32 => X"AD17DFEFA2AEAAB550051401FFA2D57FE10F7D57DE00AA842AA00007FD75FFF7",
INIT_33 => X"007BFDEAA08042AB45087FC0010557FD55FFAA843FE00F7D17FEBAA2D5574BAA",
INIT_34 => X"0000000000007BE8A005D7FEABFF002E821FF082A97555557FE8A00002E82155",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000067FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"0002074F200904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000480488024000403000000000001002A0E881108032100002000800203040",
INIT_05 => X"04092A081000411841080001000000201000012800400010001081C000402000",
INIT_06 => X"033D7880500001221021C1021800002000240249048361001100100909000222",
INIT_07 => X"9020304000220050020480152D0A142D0A8400043B45400040006810000C5901",
INIT_08 => X"0040400010880000100140024280808829029C002000000000053FA142051324",
INIT_09 => X"6008012000000000000200820888800800004000800840100020011858006442",
INIT_0A => X"000110200800840400400005C0010190070310200008B202236D080802000001",
INIT_0B => X"003000000000100C088020028102408120409120940404104C20002101004000",
INIT_0C => X"2050805210040000B0E0A0000210040000E0E0A0000190081200000000000000",
INIT_0D => X"0111300210008000B0E0A0000210008000E0E0A0000B02740421A0E5D1A02400",
INIT_0E => X"C0715C40110080A4006110510C14D18178E01200860008920106460D4501CB00",
INIT_0F => X"500002411420220080220C0093C38923240ABBC00905C33C6000400F02740412",
INIT_10 => X"9682398000120800658992F3C700C3018120000041DB011CC000090012565306",
INIT_11 => X"B7A0B1E240240A8340000200067EAA8CB65809240C09024A4AE0CA0000480083",
INIT_12 => X"00845C7DB0D0200900422ACA4B28000002002B46867DBC002A830280000800F7",
INIT_13 => X"000080020040126060008020000200000042004005800004801150A003412440",
INIT_14 => X"01088A4500008240000000802000908000800001000009A92481041000000000",
INIT_15 => X"0000000000400000000000000400000000000000000000801010000001410010",
INIT_16 => X"246810810440000090480C096420084101040000044040000000004000040000",
INIT_17 => X"4090240902409024090240902409024090240902409024090240902409024090",
INIT_18 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_19 => X"0000000000000000004090240902409024090240902409024090240902409024",
INIT_1A => X"3CF3CF3FE77DDDDD55E6D5FCF3CF3DF7CE5C8FF0F7BE9D75CF9F7DF650400280",
INIT_1B => X"FE7F3F9FCFE7F3F9FCF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"8007F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE07F",
INIT_1E => X"17DF45AAD157400007BEAAAAAAAE955555D5568A105D00000000000000000000",
INIT_1F => X"AA800AAF784020AAF7D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7D",
INIT_20 => X"0042ABEFFF8400010082EAABFF55002ABEF085155400FFD1420100055574AAA2",
INIT_21 => X"AAD540155A28028B550051574005D7FFFE105D7BD7545A284020BA0055421FF0",
INIT_22 => X"00851421FF5D7FFDEBA085168B45FF843DEBAF7843FFFFF7AABDF55A2AA97400",
INIT_23 => X"FF5504155EFAA842ABEFA280155EFFFFBC01EF08554000055002AB455D514201",
INIT_24 => X"B45557FD7410552EAAABAAA8017400AAD140000002EBFFEFA2AAA8BEFF780021",
INIT_25 => X"0000000000000000000000000000000000000000005568A1055043DEBAAAFFE8",
INIT_26 => X"F8E38E3DF45155EBD17FF6DAADB504001C71EDA82AAA0955455D556DA0049000",
INIT_27 => X"B420101C55554AAAAA480082FF84000BAEBD16DA82410A3FFD7AAA4B8E824971",
INIT_28 => X"8405092085F401D71C0A2DBC7EB80000280824ADBD7490E28BEF085157428FFD",
INIT_29 => X"BA4BDF45AAAA90410BEDF45155A28E2AB7D0051504005D71F8E004975D556DB6",
INIT_2A => X"550028B6D5D51420101C5B401EF417BFAEAA08516AB45E38E38E92EB803FFD7E",
INIT_2B => X"7A2AEAFBC7EB80071FF5500175EFB6802DBC7BE8A155EFE3FBC71FF145B42038",
INIT_2C => X"38490A3FE92BEFFEAB45417FD24385D2AAFA82B68015400AADB40000082EBFFC",
INIT_2D => X"54555557FE1000000000000000000000000000000000000000000000000556FA",
INIT_2E => X"DF45AA8428A10085568ABAA2FBD7545AAD17DFFFAAFFC200055557DE00A28015",
INIT_2F => X"A8BEF0051554AAFFFFC00105D55554BAA28400000F784020BAAAD17FE00082EB",
INIT_30 => X"568A000051575FFF78415410087BC01555D2EBFF55A284000AA08003FF55002A",
INIT_31 => X"AEA8A00A2803DF45AA843DF55AAAE82000F7FBD5545AAAEAABFF0051400105D5",
INIT_32 => X"AFBD55EF557BC20AA5D042ABFF555142000557FC01EF007FEAABA00556AB55A2",
INIT_33 => X"A2FBC0010082EBDF55A2AABDF45A284175FF5D04175FFF7803DF45FFAE955EFA",
INIT_34 => X"000000000000517FEAA082EBFE10F7FFE8B55087FC00BA552ABFE10F78415400",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000100000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"000440009282000001100000000000100220C8811080321000000228002A3000",
INIT_05 => X"04092A0010004300418800510000A6201000012A64400000145080C000422000",
INIT_06 => X"032B1800100001220001C00018821020402402080003772019001009090002AA",
INIT_07 => X"0000004000220000021840010C8912250A0400042044400040006810000C4901",
INIT_08 => X"0040400022810000058140024280A0A8190004002030C00000016F8122041320",
INIT_09 => X"E0080120000000000002C0820888008800000000800840100020011850004402",
INIT_0A => X"00013000080094000062000180010180060210200008B2022304080800000003",
INIT_0B => X"0030000000000008008020020000000000000100800000000000002500004000",
INIT_0C => X"0000000010108000000000000010108000000000000230001200000000000420",
INIT_0D => X"0000000010140000000000000010140000000000000100000040000000000000",
INIT_0E => X"0000000000000000000100008040000000000000000000020000090000000000",
INIT_0F => X"0000000030002000406000000000068409014000000000000000000100000040",
INIT_10 => X"2010000000000800000201000800000000000000400048000000000010000440",
INIT_11 => X"00184400A0000000000002000000441108800000000002008008000000000080",
INIT_12 => X"0000000242038B82800000000000000002000001000000000000000000080000",
INIT_13 => X"000080000000100000000005C04A000000400000000000000001062000000400",
INIT_14 => X"01088A4500008200000000800000100000800001000001A12480001000000000",
INIT_15 => X"4000040000000000000000000400002000020000000000801010000041400010",
INIT_16 => X"0460000004400000904808094020080000000000044040000000004000040000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000400280",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FC00000804154AA5D00001EFF78428AAA007BC2145F780000000000000000000",
INIT_1F => X"55400AA007FC2000F7D17DF45AAD157400007BEAAAAAAAE955555D5568A105D7",
INIT_20 => X"D043FFFFAAAABDEAA557BFDE00FFD140155F7FBD74AAAAD17DF45F7D1421EF00",
INIT_21 => X"F784020AAF7FFFDF45FF84000BA552ABDFEF08517DF55A2FBEAB555D556AAAA5",
INIT_22 => X"5AAFFEAB45F7843FF45082A801FF005155400FFD1420100055574AAA2AA800AA",
INIT_23 => X"AAA2D5421FF00042ABEFFF8400010082EAABFF55002ABEF087BE8ABA555168B5",
INIT_24 => X"E105D7BD7545A284020BA007FFFE10A284000AA0055401550055574005D2E800",
INIT_25 => X"0000000000000000000000000000000000000000000028B550051574005D7FFF",
INIT_26 => X"955455D556DA004971C7038140012482550E021C7EB8028A821C7BC516DFF800",
INIT_27 => X"17FF45E3DF471C70851400BA0071C5028FFD17FF6DAADB504001C71EDA82AAA0",
INIT_28 => X"FBE8B555D516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBF1D5492BED",
INIT_29 => X"C55554AAAAA480082FF84000BAEBF1FFF7DEB8000092552ABFFEF08517DF6DB6",
INIT_2A => X"087FEFA8241516DB55A2FFEAB6DEB843DF551C20801C71C5157428FFDB420101",
INIT_2B => X"5085550428412A85082BEDF401D71C0A2DBC7EB80000280824ADBD7490E28BEF",
INIT_2C => X"7D0051504005D71F8E004975D556DB68405092087FF8E00BE8A02082005F4714",
INIT_2D => X"A00557BD75EFF78000000000000000000000000000000000000000000000E2AB",
INIT_2E => X"200055557DE00A2801554555557FE100055554BA5504000105D2A80145AA842A",
INIT_2F => X"D7545AAD557410F7D57DF55AAFBD55450055420BA0055574BAF7D17DFFFAAFFC",
INIT_30 => X"ABDFFF08517FFFFF7FBEAB455D517FE00082EBDF45AA8428A10085568ABAA2FB",
INIT_31 => X"51554AAFFFFC00105D55554BAA28400000F784020BAAAD57FFEFA28402010552",
INIT_32 => X"8003FF55002AA8BEF007FFDE1000557DF45AAFBE8BEFA2803FF4555040015555",
INIT_33 => X"F7AE80000087BD55450855400BA002A95400F7FBC01555D2EBFF55A284000AA0",
INIT_34 => X"0000000000002EAABFF0051400105D5568A000051575FFF78415410087FEAA10",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000006000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"0202115002BB10080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"2FE962000017102918900948514522CE09200C0D590569398ADBF8CC1E50E480",
INIT_05 => X"5E6023002834854AE41C1E8782F508F2A15B71D412E0AFD9C2990DA56FF0B55A",
INIT_06 => X"82A803B9B9E55402000340003200220A86012D0000000480D02A7960540180A0",
INIT_07 => X"01380C40D890101DBD400901442800817C2901F400868554DE240000A80090CE",
INIT_08 => X"18A9050122004000005665510320C9C90510025A8A00000A0A048F550A440E00",
INIT_09 => X"2A8A562060410280081116C8204D016CB2CB2900080082795804112890000001",
INIT_0A => X"4052E400008176802200020025699200140001A15000017F0051D0F837324E00",
INIT_0B => X"5514554485D000000124002400000000000001004010A8812831605DA0000A05",
INIT_0C => X"708E2CB5320018CAC99BA0A3B9320018CAAAADA0C343F1AC1B01040A00202489",
INIT_0D => X"E7A3EE59320018CAC99BA0ACB9320018CAAAADA0CC421CA003B694B68018FAAA",
INIT_0E => X"24352AB2449A3FF2FA04E5E09B128834ADB1443A1891E4A928C29020E6A8524C",
INIT_0F => X"714C902375B801324301AB0067622E5E5404B2A5A40B1E6644AF0F021EA003AC",
INIT_10 => X"1216F50A8C241815FEB6A9158863F638FB60ED838E890B703C6260D8E3A21275",
INIT_11 => X"555E4C15F11133D171727A2550EE2F1BA0064F70DBDB1C74424E91E1C194C71D",
INIT_12 => X"ACCC59432A2B2D001F803471A9A960E57245FDF9D364DBD9435A6D45C9E81BED",
INIT_13 => X"0012CAC00006B0800000038814B72AB01508150013F162119014204373517700",
INIT_14 => X"002912300208092B940192D1000000000000A8A5AA80018120E0006600000000",
INIT_15 => X"1100011000110001100011000108000880008000520228080108039501200848",
INIT_16 => X"012000081500008A422150884081AC9000010003561180063DB4F61100011000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"28A28A3D2DE5F87963445469E79E7853D44C690DA64C1C69818768A360400000",
INIT_1B => X"F4FA3D3E8F4FA3D3E9A29A29A29A29A29A29A29A29A29A29A29A29A28A28A28A",
INIT_1C => X"000FA7D3E9F4FA7D1E8F47A3D1E8F47A3D1E8F4FA7D3E9F4FA7D3E9F4FA7D3E8",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"43FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE005500000000000000000000",
INIT_1F => X"80020005D2A95410FFFFC00000804154AA5D00001EFF78428AAA007BC2145F78",
INIT_20 => X"AD157400007BEAAAAAAAE955555D5568A105D2E974BAF7FBEAB45FFFFC00BAF7",
INIT_21 => X"007FC2000F78000010552E800AA002E821FFA2AAAAA00000417555FFD17DF45A",
INIT_22 => X"A08043FEBA5D55575FFF7AABFE00557BD74AAAAD17DF45F7D1421EF0055400AA",
INIT_23 => X"10FFD56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7AABDF55F7AE820A",
INIT_24 => X"FEF08517DF55A2FBEAB555D04154BAA2FBE8B55FFFFD55FF557FC2000FF80154",
INIT_25 => X"0000000000000000000000000000000000000000007FFDF45FF84000BA552ABD",
INIT_26 => X"28A821C7BC516DFF8438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE1049000",
INIT_27 => X"BE8B55FFF1C70BAF78A000005D2097438FFF1C7038140012482550E021C7EB80",
INIT_28 => X"0E1757DEBD17FF6DAADB504001C71EDA82AAA0955455D556DA00492490492F7F",
INIT_29 => X"3DF471C70851400BA0071C5028FF84020285D2085092002A801FFB6AAA8A1008",
INIT_2A => X"EBA4BAF6DE3AA8709208043FEBA555B555FFE3AABFE005D71D5492BED17FF45E",
INIT_2B => X"7557BC0028E38412428EBD16DA82410A3FFD7AAA4B8E824971F8E38E3DF45155",
INIT_2C => X"7DEB8000092552ABFFEF08517DF6DB6FBE8B555D04124BAB6FBE8B45E3FBD55D",
INIT_2D => X"55555003DE000000000000000000000000000000000000000000000000071FFF",
INIT_2E => X"00105D2A80145AA842AA00557BD75EFF78428B55AAD168B55F7FFFDFEFFFAA95",
INIT_2F => X"7FE10000000010F7FBEAB45FFD1554AAFFAE820105500154AAF7D5554BA55040",
INIT_30 => X"E801EFF7AEA8A10002E955FFA2D17DFFFAAFFC200055557DE00A280155455555",
INIT_31 => X"5557410F7D57DF55AAFBD55450055420BA0055574BAF784000BA5D0017410082",
INIT_32 => X"85568ABAA2FBD7545AA802ABEFA2AA9541000003DEBA557BD75EFA2AEBDE105D",
INIT_33 => X"FFFBEAB45AAFFD55555D7FC20AAA280000AAAAD17FE00082EBDF45AA8428A100",
INIT_34 => X"000000000000557FFEFA28402010552ABDFFF08517FFFFF7FBEAB455D04020AA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000002000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"5295B6957FCBE0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"6DE90201BF90102103AF158E805428249851BFB2C106592088DBF8400A5055C2",
INIT_05 => X"3824BD7F80148D9E07100A8201ED01C1A19B68F40A807ED9C18114956FF081DB",
INIT_06 => X"ED08CA6A8F033DD800000000050716BE9F57F8AC000807DFD999E0E5E1818B1B",
INIT_07 => X"00150886481240FE05A109228E2C0891D772A6F40045B8CF30E085DD2ED57D4E",
INIT_08 => X"72637FDF23800005981C0338190549C904182B6113870022000488C08B46268A",
INIT_09 => X"3E7437823DF78CDB6CA60E0E28EFFE2061872F80C1684A80C8604085F0074D3B",
INIT_0A => X"F5B4FFBD2FAD7FE653C36A1FF33E0E001E000B3A5DAADAFDDA5DA79350CFB801",
INIT_0B => X"CFE833C5C3D00018006C681700000000000000020012E9E10A31EB5FF9296A67",
INIT_0C => X"0D5ECE542A6FEEB2533EA160782A6FEEB2333EA16031F2BD47BDA2CA5D8164FC",
INIT_0D => X"282400F82A6FEEB2533EA160782A6FEEB2333EA160391BEFF2C32FB695F91911",
INIT_0E => X"573FAD5A86840354D1706FFFA3EF6E24B6D18C0D06638A207CFDE1F7DDAD76D5",
INIT_0F => X"FE4ACA4D77FAAB77CE3AF3EE78F58DB737E6E43E59AFE4A59B57679D19EFF2C7",
INIT_10 => X"ADB55572CA52606DFED6CA55334C04C04FF7D7A0ABD6DAAAB96529382B74E4E1",
INIT_11 => X"F9956EAA1A184045D5D7A870D2F5A5D7522D1281017F056E9C9C3FC95949C157",
INIT_12 => X"1F432EA58949D5B5C85F97871876F7D7E859FDEB974F486905001FDF5FA0D719",
INIT_13 => X"DEF20670021EE341036BF368128419FB5560158015177F916A039EF41FDB34A9",
INIT_14 => X"00633F1D0A7CC9AE7A08BFF0001D35682AC0CE8FCCC200A59BDD2FFE3F3EC7C7",
INIT_15 => X"FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A7800617112E46F05D02DD814102F8",
INIT_16 => X"05F08000179C16DECF67F08BC02F9086000D9E8A3F06ABD73DBCF4FBCF4FBCF4",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"34D34D48C4986868DC800181D75D7445F009EDCC4052E92E0204114F981800C0",
INIT_1B => X"1A8D468341A8D46834D35D74D34D35D74D35D74D34D35D74D35D74D34D34D34D",
INIT_1C => X"0008D46A351A8D46A351A8D46A351A8D46A351A0D068341A0D068341A0D06834",
INIT_1D => X"0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"43FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF5500000000000000000000",
INIT_1F => X"8028A00F7843FEBA55043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE00550",
INIT_20 => X"804154AA5D00001EFF78428AAA007BC2145F7D568B45000002010552EBDF45A2",
INIT_21 => X"5D2A95410FFAE800105D2A95410002A95410AAAEBFF55AAFFC00BAF7FFC00000",
INIT_22 => X"FFFD57DE00F7AE800AAAAAABDFEF5D2E974BAF7FBEAB45FFFFC00BAF78002000",
INIT_23 => X"AA5D517DF45AAD157400007BEAAAAAAAE955555D5568A105D7FFFFEFA2D568BF",
INIT_24 => X"1FFA2AAAAA00000417555FF8028B55082A974105D003FF55F7802AAAAAAD168A",
INIT_25 => X"0000000000000000000000000000000000000000000000010552E800AA002E82",
INIT_26 => X"955C71C043FE10490A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD749000",
INIT_27 => X"E050384124BFF7DB68A28A38F7803DE82490438FC7E3F1EAB55B6DF6DBFFF7AA",
INIT_28 => X"F5C70BAFFF1C7038140012482550E021C7EB8028A821C7BC516DFFDF68B551C0",
INIT_29 => X"FF1C70BAF78A000005D2097438FFAA85000492495428082E95400AAA0BDF7DB6",
INIT_2A => X"497FFAFFFB6D56FBFFEBDB78E38F7AA800BAB6AEBDFD75D2490492F7FBE8B55F",
INIT_2B => X"DEB8028AAAB6D16FA8249517FF6DAADB504001C71EDA82AAA0955455D556DA00",
INIT_2C => X"285D2085092002A801FFB6AAA8A10080E1757DEB8A2DB5514249243841003FF6",
INIT_2D => X"0BAF7FFFDF550000000000000000000000000000000000000000000000004020",
INIT_2E => X"8B55F7FFFDFEFFFAA9555555003DE00002ABFFEFF7FBFDFFFAAD168B55AA8000",
INIT_2F => X"D75EFF7FBEAB45552E954BA08003DFFFFFAAA8AAAF7843FE10000428B55AAD16",
INIT_30 => X"E95410AA843FFFFF7D5554BAF7D5554BA5504000105D2A80145AA842AA00557B",
INIT_31 => X"0000010F7FBEAB45FFD1554AAFFAE820105500154AAF7AE974000800154AA002",
INIT_32 => X"2801554555557FE10007FEABEFFFD57FFEFAAFFE8ABAFFAA820BAF7AEBFF5555",
INIT_33 => X"5500020AA08003DFFFA28028AAAF7D17DE0000517DFFFAAFFC200055557DE00A",
INIT_34 => X"00000000000004000BA5D0017410082E801EFF7AEA8A10002E955FFA2AABFF45",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000067FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"080BA868803F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"42016B0C401F58495C900A4859552A611D9A640F5903B2388004004C08A06008",
INIT_05 => X"16226B107811422A641C08038040007060E0032801E0202000991B708280B501",
INIT_06 => X"120886B3B8E0FC86142B4142B0000000011114D3058240240907F82000000000",
INIT_07 => X"006880802102401015610A02C4005000EA019D002482043FCF1C8090C02800C0",
INIT_08 => X"11018020D40A5004003260F9810541494D403D9B98810A0002C601000054B94A",
INIT_09 => X"022E0C6070000504102805C820C8016C30C250080C0182183804012A0A102200",
INIT_0A => X"084001E000108010230495A800FD865421432121804021C20452880C2D100000",
INIT_0B => X"3F140FC2060014250B9080008306C18360C1B0609C05013065CC042004040808",
INIT_0C => X"DF7C728582081483ACC15F9C3982081483CCC15F9CBA45505640000A40201900",
INIT_0D => X"DFEBFBF982081483ACC15F9F3982081483CCC15F9FB1962FCB69E08AAAEAEBCD",
INIT_0E => X"CAA02FE3F8E7F5E3AC3620805298B15A3FEBF1CFFF7670ACC3811A28AB57523C",
INIT_0F => X"01BD67DC4041D4CF03138DD865103EFEEAC9002BF05800D875E63CC9962FCB52",
INIT_10 => X"0016EA8DB7BFE25208E8F46A228BF8A757F1B72A8A800B7546DB9F1CA320037F",
INIT_11 => X"81A8A29509EAAE7FD3B749471C48F8A45981CCFAFDBF9464006FD037AEFAE515",
INIT_12 => X"EFF5778802A3AF8E8FB0440CE78773B709641256EC844B8AF92FD7CEDC24A9E1",
INIT_13 => X"0003C1C284601C2864000080113307E4800297D086E00036D2440E0880AAD62B",
INIT_14 => X"C44C92A88DCC2211E44174112840880000060D7030C30B885200D27400400808",
INIT_15 => X"0030800308003080030800308001840018400400602A01880980037109700C04",
INIT_16 => X"6808348340000020301805002D008CD943626111C0D95C20C2030A0030800308",
INIT_17 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B0",
INIT_18 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_19 => X"00000000000000000041B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_1A => X"1451451223059150A2EFB05C104104B3CEB80EE173C2300FCA8B7DF160000000",
INIT_1B => X"4AA552A954A25128955545145145155555545145145155555545145145145145",
INIT_1C => X"00025128944A25128944A25128944A25128944A25128944A25128944A2512894",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"43FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA0000000000000000000000",
INIT_1F => X"8400145AA801741000043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF550",
INIT_20 => X"7FBE8B45AAD568BFFFFAA975FF00003FE0055043FFFFFFFFFDFEFA2D56AB45AA",
INIT_21 => X"F7843FEBA55557FFEFA2D168B55AAFBFFFFFFF80021EF0855421EF00043FFFFF",
INIT_22 => X"A5D2A82155F7AEBFEBAFFD56AA00A2D568B45000002010552EBDF45A28028A00",
INIT_23 => X"BAA2FFC00000804154AA5D00001EFF78428AAA007BC2145F7D5400000004020A",
INIT_24 => X"410AAAEBFF55AAFFC00BAF7AE80010082E954BA0004174AAAA8428B45082ABFE",
INIT_25 => X"0000000000000000000000000000000000000000002E800105D2A95410002A95",
INIT_26 => X"00038F7DB6FBD7490E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA55041549214000",
INIT_27 => X"1F8FD7AAD16FB6DBE8E00155BE8015410140A3FFFFFFFFFDFEFE3F5FAF45AA80",
INIT_28 => X"5B471C7140438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE1049043FFEFE3F",
INIT_29 => X"124BFF7DB68A28A38F7803DE82495B78FC7AAD56FB6DBEF1FAFD7E384001EF14",
INIT_2A => X"FFD1420381C0A02082492A85155E3A4BDE92FFD56FA28B6DF68B551C0E050384",
INIT_2B => X"ABE8E28B7D1420BDEAAA2F1C7038140012482550E021C7EB8028A821C7BC516D",
INIT_2C => X"00492495428082E95400AAA0BDF7DB6F5C70BAFFAE870280024904BA1400174A",
INIT_2D => X"4BA550415410550000000000000000000000000000000000000000000002A850",
INIT_2E => X"DFFFAAD168B55AA80000BAF7FFFDF55002ABFFFFFFFFFFFEFF7FBFDFFFF7AA97",
INIT_2F => X"3DE0000043DFEFA2D56AB45AAD57DFEFF7AA82155F78015400552ABFFEFF7FBF",
INIT_30 => X"568B55A280021EF557FD7555550428B55AAD168B55F7FFFDFEFFFAA955555500",
INIT_31 => X"FBEAB45552E954BA08003DFFFFFAAA8AAAF7843FE10007FEAB55A2D17FFEFFFD",
INIT_32 => X"A842AA00557BD75EFF7D1400AA5D2A82000002A95545A2843FE00F7D17FEAAF7",
INIT_33 => X"0004020AA5D04154BAF7AEA8BEF55003DEAAA2D5554BA5504000105D2A80145A",
INIT_34 => X"0000000000002E974000800154AA002E95410AA843FFFFF7D5554BAF7AE974BA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000002000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000010228001000000000000000000024001620280000000000354200004008",
INIT_04 => X"00016200001310090090004840004152C7208802590000388000004C08006000",
INIT_05 => X"1621008008100002641C0803804000702000000000E02000009900000000B100",
INIT_06 => X"00A0010210200C00000000000000000000000080000000000000D82000000000",
INIT_07 => X"010084C00D267001B880080700285020020AC988200228024004804050089011",
INIT_08 => X"0E0E00000000000000106009872048400C4000010D000008000204150A00815A",
INIT_09 => X"022A040000000000000004C80000002C30C20000000002180800580000000000",
INIT_0A => X"0007600000000000000000080025860000000080A00020602040800000000000",
INIT_0B => X"031400C002000000000000000000000000000000000000000000000000000084",
INIT_0C => X"28DC0D385598035D0008A003B05598035D0008A0034078104B41A41000000000",
INIT_0D => X"041124505598035D0008A000B05598035D0008A0004263C0343EDD4140040422",
INIT_0E => X"B740500401180DE053A98F6ECC739D8140040231068187C39F5A4F985C008902",
INIT_0F => X"000010227848D4303807FC8CC5508AEAED1BFBD406451B02000E033263C0343C",
INIT_10 => X"D6480000000018A700FCF980CC300318A2420851546B2400000040D8549B5800",
INIT_11 => X"81C21140E40511802208D6B30C48F8A8A452210402120A936B0000000004C2A8",
INIT_12 => X"F9E9410006362A2B6424287B08286208D6B1427ED430B41402D0250823597001",
INIT_13 => X"0002C040000000000000000010030060009C000018440021011821B35254E99A",
INIT_14 => X"000040002000044000000000000000000002F0001F00002024B2000200000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"00000000000000000000000000008C8000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C30C30D0A208C4DC822EC1534D34C01FA3F0C7010C6600A0200441920000000",
INIT_1B => X"26130984C26130984C30C30C30D34C30C30C30C30D34C30C30C30C30C30C30C3",
INIT_1C => X"000130984C26130984C26130984C26130984C26130984C26130984C261309A4D",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D00000000000000000000",
INIT_1F => X"AA974BA5D517FFFF08043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA007",
INIT_20 => X"FFFFFFFFF7FBFDF55A28402000F7D56ABFF557BFFFFFFFFFFFFFFFFFBFDFEFFF",
INIT_21 => X"AA8017410007BFFFFFFFFFFFFEFF7D16AB45AA8002000F7D5575455D043FFFFF",
INIT_22 => X"5AAD568B55F7AE955FFAA840201008043FFFFFFFFFDFEFA2D56AB45AA8400145",
INIT_23 => X"FF5D043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE00557BFFFFFFFFBFDF4",
INIT_24 => X"FFFFF80021EF0855421EF002ABFFEFF7D168B55AAD17FFEFF7AE975FF00557FF",
INIT_25 => X"000000000000000000000000000000000000000000557FFEFA2D168B55AAFBFF",
INIT_26 => X"954AA5504154921471FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA55000008255000",
INIT_27 => X"FFFFEFF7FBFAFD7E3A4954BA555B7AFC7080E3FFFFFFFFFFFFFFFFBFDFEFFFAE",
INIT_28 => X"DF52545550A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD74975FFFFFFFF",
INIT_29 => X"AD16FB6DBE8E00155BE8015410147FFFFFFF7FBF8FC7EBD568B55A28000000FF",
INIT_2A => X"497BFDFC7E3F1FAF55A2DB6FB7DF7AE955C7BE800000008043FFEFE3F1F8FD7A",
INIT_2B => X"7EBA0955FF145B7AFC7410438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10",
INIT_2C => X"C7AAD56FB6DBEF1FAFD7E384001EF145B471C71424B8FC7E3D56AB6DB6DF7AFC",
INIT_2D => X"4AA550002000550000000000000000000000000000000000000000000005B78F",
INIT_2E => X"FFEFF7FBFDFFFF7AA974BA55041541055517FFFFFFFFFFFFFFFFFFFFEFF7AA97",
INIT_2F => X"FDF5500517FFFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB45002ABFFFFFFFFF",
INIT_30 => X"56AB55A28002000F7FFC2155552ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FF",
INIT_31 => X"043DFEFA2D56AB45AAD57DFEFF7AA82155F78015400557BFDFEFF7FBEAB55A2D",
INIT_32 => X"FAA9555555003DE00007FFDF45AAD568B45AAFBFFFFFFFAA95545F7840201000",
INIT_33 => X"AAD16ABFFFFFBEAB45A280155EF557FE8B55000428B55AAD168B55F7FFFDFEFF",
INIT_34 => X"0000000000007FEAB55A2D17FFEFFFD568B55A280021EF557FD755555042AB55",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000004000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"0001E6000053300B00D0005800000000000000407B0004BB830004DC3D01E000",
INIT_05 => X"FEE0000008720043EC3C3D0F87FA19F7E0201C409BE1F10623BB000A100CF300",
INIT_06 => X"00200006102FFC8E0007C00078008000171175A200096404D97FFBE4744200AA",
INIT_07 => X"000000482491301000010001DC00000000000000004203FE4005800000008030",
INIT_08 => X"40800020E2008000027FEFF946058180010429000001080AAA010F8000000000",
INIT_09 => X"03EAFE400000120000913FD80000003DF7DE0080010047FBF8000000000800C5",
INIT_0A => X"0800000080000010000400080FFDBE0000004000000100000100506002204610",
INIT_0B => X"FF14FFC00600000000801020000000000000010240001721214E000004000000",
INIT_0C => X"A70C0008020000200000000F30020000200000000F3008001E00000000001803",
INIT_0D => X"004A58F0020000200000000F30020000200000000F3040200000020000000026",
INIT_0E => X"000000000019B140000800800000020000000030B86000400080000200000000",
INIT_0F => X"000014AC08000000508001030A0A4001000000000002183E61E6000040200001",
INIT_10 => X"0000000000A56000090100000000001F86C00010080000000000525801000000",
INIT_11 => X"0600000000001716800000803102020000000002BC360020000000000292C010",
INIT_12 => X"06049CDF70C08040100000706707600000801000000000000057450000100106",
INIT_13 => X"000ADFC011001C81080001101F977FE008000000000000400400400020000805",
INIT_14 => X"0000000000000000000000020020029000000000000000020000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000002000200000000",
INIT_16 => X"0080800801810100000000000093ED8000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000401",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"18618640C49821201C0001A1E79E79A4B0038200010089054C1A0104D2040020",
INIT_1B => X"0C86432190C86432196596596596596596596596596596596596596586186186",
INIT_1C => X"00086432190C86432190C86432190C86432190C86432190C86432190C8643219",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA5504020100800000000000000000000",
INIT_1F => X"AA974AA550002000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7",
INIT_20 => X"FFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFFFFFFFFF7",
INIT_21 => X"5D517FFFF087FFFFFFFFFFFFFFFFFFFFDFEFFFAE974AA5D003FE005D043FFFFF",
INIT_22 => X"FF7FBFDFFFAA84000105D556AB55557BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA",
INIT_23 => X"EF08043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55003FFFFFFFFFFFF",
INIT_24 => X"B45AA8002000F7D5575455D2EBFFFFFFFFFFFEFF7FBEAB55A28000010F7D16AB",
INIT_25 => X"0000000000000000000000000000000000000000007BFFFFFFFFFFFFEFF7D16A",
INIT_26 => X"954BA550000082557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA55040002800000",
INIT_27 => X"FFFFFFFFFFFDFEFF7AE974BA5500050380071FFFFFFFFFFFFFFFFFFFFFFFF7AA",
INIT_28 => X"0038E285D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA55041549214043FFFFFFF",
INIT_29 => X"7FBFAFD7E3A4954BA555B7AFC70871FFFFFFFFFFFFFFF7FBFDFFFFFAA974BA55",
INIT_2A => X"490E3FFFFFFFFFDFEFF7F1FAFC7A28002028555F6FB7D5D75FFFFFFFFFFFFEFF",
INIT_2B => X"5A28402010FFDB6ABEF140A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7",
INIT_2C => X"FFF7FBF8FC7EBD568B55A28000000FFDF525455524BFFFFFFFBFDFC7E3F5E8B4",
INIT_2D => X"4AA5504000BA080000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFEFF7AA974AA550002000557FFFFFFFFFFFFFFFFFFFFFFFFFFAE95",
INIT_2F => X"1541055043FFFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08517FFFFFFFFF",
INIT_30 => X"FFFFEFF7AE974AA550028AAA5D2ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA5504",
INIT_31 => X"517FFFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB4500557FFFFFFFFFDFEFF7F",
INIT_32 => X"A80000BAF7FFFDF55002EBFFFFF7FBFDFEFFFD568B55A284020BA557FFFFFF5D",
INIT_33 => X"F7FBFFF55A2D16AB45AA8402000F7FBEABEF5D2ABFFEFF7FBFDFFFAAD168B55A",
INIT_34 => X"0000000000007BFDFEFF7FBEAB55A2D56AB55A28002000F7FFC215555043DFEF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"1094EC681244819000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"0001E6000053300F01D4587800446194F49020107F0012BBC00202DC3823EA82",
INIT_05 => X"FFF201B228704123FC3C381F87C03DFFF012412A9FE1E01013BF09404050F300",
INIT_06 => X"100B3096F43FFF002004020044041084CB01AD0000037617027FFFE050000080",
INIT_07 => X"A12034043C802A821D41412001A0040950AB60014114C3FE4187A009A663A680",
INIT_08 => X"7F40002C01004000047EFFF811A46968004060629A0002208A00000068113205",
INIT_09 => X"E3EBFE0A812D8D5B742D3FF84056383FF7DE0880042107BFF9C45B85101C49A3",
INIT_0A => X"02804A08221890004806C0310FFDFE00040009814C089202225412115414601D",
INIT_0B => X"FF56FFC0281280080180B2948004400220011100841200D001000624000100C0",
INIT_0C => X"50025360694101816002D41A4068C101815004D8158809C86065941840B1014F",
INIT_0D => X"82418A0068C101816002D41A40694101815004D815810D42E04A08A80098C024",
INIT_0E => X"1A300012682960828F05C96A001B029010134160C8125B0B271802242880A044",
INIT_0F => X"49F115100920C54E8EA256ECF078BA081C10080E05C0B06AA8B12CFD0D42E044",
INIT_10 => X"5144104F30A8801406D00290006280320100010362A8A20826A88660D86B2020",
INIT_11 => X"8010602011819E290048A2118EC8140C08064802C0081B0D64040936443306C5",
INIT_12 => X"C322A4C40A0300600C0A80509F418008804581BA0038005A706680012280506A",
INIT_13 => X"18DBFFC000120080002341881F3FFFF80DCC158092C044600466208CC5091011",
INIT_14 => X"806520398C6021569249C4B3007127080806FF917FC30010107688862A28C545",
INIT_15 => X"9228D9228D9228D9228D9228D99146C9146C84006309044081A001B188300E20",
INIT_16 => X"0448008004000000E07008010003EF80022A51904595123203040D9228D9228D",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_19 => X"0000000000000000004010040100401004010040100401004010040100401004",
INIT_1A => X"7DF7DF7FEFFDFDFFFBE7F3FCF3CF3FFF6EFF7FFDF7FF3EFC1FBFFDF7E0000000",
INIT_1B => X"FEFF7FBFDFEFF7FBFDF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF",
INIT_1C => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFD",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D00020000800000000000000000000",
INIT_1F => X"AE954AA5D00020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"55000200000003FFFFFFFFFFFFFFFFFFFFFFF7AA974BA5D0402000557BFFFFFF",
INIT_22 => X"FFFFFFFFEFF7AE974BA5D00174BA00003FFFFFFFFFFFFFFFFFFFFFFF7AA974AA",
INIT_23 => X"BA5D043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFF",
INIT_24 => X"FEFFFAE974AA5D003FE005D2EBFFFFFFFFFFFFFFFFFFDFEFF7AE954AA5500174",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFD",
INIT_26 => X"974AA550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000001000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"04050005571FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082557BFFFFFFFF",
INIT_29 => X"FFFFDFEFF7AE974BA55000503800003FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D",
INIT_2A => X"140E3FFFFFFFFFFFFFFFFFFDFEFF7AE954BA5D00154AA00043FFFFFFFFFFFFFF",
INIT_2B => X"FFFAA974BA5D00104925D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492",
INIT_2C => X"FFFFFFFFFFFF7FBFDFFFFFAA974BA550038E285D2ABFFFFFFFFFFFFFFFFBFDFE",
INIT_2D => X"4BA5D00000100000000000000000000000000000000000000000000000071FFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02000557BFFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7FFFFFFFFFFF",
INIT_30 => X"BFDFEFF7AE954AA5D041740055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5500",
INIT_31 => X"043FFFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08043FFFFFFFFFFFFFFFF",
INIT_32 => X"7AA974BA550415410552ABFFFFFFFFFFFFFF7FBFDFFFFFAA974AA5D00174BA08",
INIT_33 => X"FFFFFDFEFF7FBFFFFFF7AE954BA5D0000010552ABFFFFFFFFFFFEFF7FBFDFFFF",
INIT_34 => X"000000000000557FFFFFFFFFDFEFF7FFFFFEFF7AE974AA550028AAA5D2EBFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"8632CA211E4491D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"24B000808800040439245B221373581F97B0A8D1040F92000F42000047A00E58",
INIT_05 => X"011B2BBA308F023810004700083E220811E9BF2844021B1004045E4249500449",
INIT_06 => X"EF018980A51003AA0200C020088E16A85235722940A817251100040D6D0702A2",
INIT_07 => X"24E8145C9ECAB0D247B013B405EAD525FAE48FC2060B880081A26DCD4047EFF9",
INIT_08 => X"0050482D0141C0055280100751096B6A40D6F86723E510AA2004803D3275EB20",
INIT_09 => X"20110204804818CD280100207246A8020000AC0283002004051507A5411C0DA0",
INIT_0A => X"4E506A2C6898B2950AA6D635B00041C23020131A80CFDFF3FE509A907C556828",
INIT_0B => X"002200050F60E220A06880D2A14050A028501428054278142151262CA5034385",
INIT_0C => X"F06273612B3482C0C0078E1F412B1582C090078E1F840A2B0114020104022460",
INIT_0D => X"C2C0DB012B1582C0C0078E1F412B3482C090078E1F891C239F8908003099C1AC",
INIT_0E => X"0828041BA859F213AFC14AA380430060181BA1B0FD16770236A4091621C08055",
INIT_0F => X"095337B08AA600CA88B143AB11880C280600101F09C030AB28B03C111C239F87",
INIT_10 => X"3096004B61BD8068B92400D0004E30368910E8822A984B0025B0DE6089462660",
INIT_11 => X"F07830001AC2173B00E162563454C40804055412D4481128C4CC012A66F30455",
INIT_12 => X"BF006850840180A00E1C81900C4190E160589C48082C006A9057CA4385809520",
INIT_13 => X"39C020004416B105036B4180C000800C8C00460848952220592745AC11A544B1",
INIT_14 => X"103D2A512C6A8C4F0008AA800470370000A0004D0000002126F30C902A29C545",
INIT_15 => X"C2A81C2A81C2A81C2A81C2A81C9540E1540E001400006100003202D040050220",
INIT_16 => X"45E22022365034A8EA754008004C0214202C50013456520CA09281C2A81C2A81",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"0040100401004010040100401004010040100401004411044110441104411044",
INIT_19 => X"0000000003FFFFFFFF9004010040100401004010040100401004010040100401",
INIT_1A => X"3CF3CF7FE7FDFD7DF7EFFDDDF7DF7DF7DEFE8FF1F7DEBD6FCD9F7DF7D0512289",
INIT_1B => X"FE7F3F9FCFE7F3F9FCF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"0007F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04000000000000000000000000000",
INIT_1F => X"AE974BA550000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D00020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00000AA007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAA954BA5504000AA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA",
INIT_23 => X"BA5D7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFF",
INIT_24 => X"FFFF7AA974BA5D040200055517FFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500000",
INIT_25 => X"000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040200008000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"00020BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D",
INIT_2A => X"5571FFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5504020AA5D7BFFFFFFFFFFFFFFF",
INIT_2B => X"FF7AA974AA5D00070925D71FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082",
INIT_2C => X"FFFFFFFFFFFFFFFFFFEFF7AA974AA5D040500055517FFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D040200008000000000000000000000000000000000000000000000003FF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAA954AA5D00020AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504",
INIT_31 => X"7BFFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7BFFFFFFFFFFFFFFFFF",
INIT_32 => X"7AA974AA55000200055517FFFFFFFFFFFFFFFFFFFFEFF7AA974BA5504020BA55",
INIT_33 => X"FFFFFFFFFFFFFFDFEFF7AE974AA5D00154105D517FFFFFFFFFFFFFFFFFFFFEFF",
INIT_34 => X"000000000000043FFFFFFFFFFFFFFFFBFDFEFF7AE954AA5D041740055557FFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"5886C0201A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"0005EE040057700F40D08078500000D9218020407F0000BB8018A2FC380BEAC2",
INIT_05 => X"FFE0419028700023FCBC385F87C0BFFFE0124002FFE1E0C517FF09111212F300",
INIT_06 => X"DF0AF116D03FFC96102081020000020489019C4304802412027FFFE000000000",
INIT_07 => X"B710000001160A003475C8100123400E20E1F40F439647FF4807E189A477EF81",
INIT_08 => X"7F0F94801008000007FEFFFB110140695812CC4188D58A0AAA10803448D0844F",
INIT_09 => X"C3EBFD4201258112D4487FF8001010FFF7DE4000000003BFF8C2581808002001",
INIT_0A => X"0801000C024000004A9400000FFDFF50010103134CAFDF03BA18000F39900037",
INIT_0B => X"FF57FFC02812F00429DC92C40002000100008000105400C00400100000A01800",
INIT_0C => X"424202A1CAF13F214001521001CBF03F21100152100801C17E61841950B1C10F",
INIT_0D => X"420B8001CBF03F214001521001CAF13F2110015210088528E00E02C8200A430A",
INIT_0E => X"12480202C86040902AC60BACDF0E02D02001C1C044006D0C94FB94320880603C",
INIT_0F => X"09B00300010AF5052419D196441902801430182800A018D9CA8000648528E00D",
INIT_10 => X"C140004D101808458A5602E000892029110445C19960A00026880C0067390000",
INIT_11 => X"4040301009408021144CB042F880100C0601844068880CE72000013600600332",
INIT_12 => X"EE38A1F80E02120018390320F050144CB241D0B9023402085020825132C8CB5B",
INIT_13 => X"001BFFC200400020224000405F7FFFE0008E17C0D240406519400500840A9524",
INIT_14 => X"907120AC810033149249C433200180082A06FF907FC308181204800600000000",
INIT_15 => X"1010C1010C1010C1010C1010C10086080860840063090442A18001B188300C48",
INIT_16 => X"2000100100000000000004002403EFC10302219A41C1443243050C1010C1010C",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_19 => X"0000000000000000000080200802008020080200802008020080200802008020",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"550000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974AA550400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"00087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE954AA5D00000AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA5504020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA55",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400010087FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE954AA5D0402038007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE954AA5D00020BA087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"00010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D00",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA55040001000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAA954AA5D04000AA087FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D00020AA007BFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"0000745C200801000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"0001E6000053300F00D0007810042140C00000407F0000BB800000DC3801EA00",
INIT_05 => X"FFE0000008700003FC3C380F87C019FFE01240009BE1E00003BF00000000F300",
INIT_06 => X"DC8C3006103FFC0000000000000000048900880100800012027FFFE000000000",
INIT_07 => X"0061200009B24B043980021000810284204A8001401643FE4007E5501AA00000",
INIT_08 => X"7F00000000000000007EFFFB11A56940581280031D61420000B080102040BC5B",
INIT_09 => X"C3EBFC020125811254083FF80000003FF7DE0000000003BFF800580000000001",
INIT_0A => X"0580000000000000000000000FFDFF4000000AA0354000019C40000128000011",
INIT_0B => X"FF56FFC000104000000010440000000000000000001000C00000000000000240",
INIT_0C => X"48C0804012500021B00880108012500021E00880104809C1666594584031010F",
INIT_0D => X"0501840012500021B00880108012500021E0088010492064206100E810842000",
INIT_0E => X"0270040410004C840041A0D8005410903804100144800803419043064900C002",
INIT_0F => X"400041020902F60002260D65B361BAA1041018140F02C0000809408D20642053",
INIT_10 => X"D0021800020818B06D9802F00030C02060110002C9E8010C00010480B35A0300",
INIT_11 => X"90203020042108603100061516EE800C060228204300166B4060080008240593",
INIT_12 => X"14AE4C7C02000040206602C10B48110006143B62023C00142800B04400095DFF",
INIT_13 => X"001BFFC000000000000000001F17FFE000DC1180C78044000440292083010402",
INIT_14 => X"814080008000010012414433000100080806FD107FC300000000000600000000",
INIT_15 => X"1000C1000C1000C1000C1000C100060800608400630104408180012188300C00",
INIT_16 => X"0000000000000000000000000003EF80020201904181003003000C1000C1000C",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"3DF3DF64C7986120B42BB99575D75FFD2AF6E7CC1132CD73DF3A441990000000",
INIT_1B => X"1E0F0783C1E0F0783DF7DF7DF7CF3CF3CF3CF3CF3DF7DF7DF7DF7DF7DF3DF3DF",
INIT_1C => X"0000F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100800000000000000000000",
INIT_1F => X"AE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"00007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D00020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010080000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000001008",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA550000010087FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002010087FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00004000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"4909E6093253306F82D0007C80000000080E01007F8020BBC00040DC3801EA00",
INIT_05 => X"FFE0000008704503FE3C380F87C019FFF01241009BE1E00203BF80800000F392",
INIT_06 => X"CC083006103FFF9E2086C2086E006604C9019D03108B7412027FFFE070400880",
INIT_07 => X"0000004024057000000100000000000000000001401643FE4007C00000000000",
INIT_08 => X"7F00000801404000007EFFFF40010000401408000045000000A0801000408000",
INIT_09 => X"C3EBFF4A7DF795965C6D3FFC0020003FF7DF01880C618FBFFDD75E0010004043",
INIT_0A => X"0000000000000000009400000FFDFFC006020000000000019804000028000191",
INIT_0B => X"FF56FFC02812E0182000F2C48304418220C11160845004D04820000000000000",
INIT_0C => X"0800800002400001000800000002400001000800000801C0786184185031810F",
INIT_0D => X"0400000002400001000800000002400001000800000000202000000800000000",
INIT_0E => X"0200000000000404000000880000001000000001000000000090000008000000",
INIT_0F => X"000040000100C600800001040000040009100000000200200000400000202000",
INIT_10 => X"4000000002000000081001000000000040010000082000000001000001080000",
INIT_11 => X"0000400080000040010000001080001008000000010000210000000008000010",
INIT_12 => X"0420000000030280000000010000010000001020000000000000100400000108",
INIT_13 => X"001BFFE0120012C1400080291F17FFF0018C11808200400000400000C2000000",
INIT_14 => X"80400000800001001243443B000100880806FD107FC301800000000600000000",
INIT_15 => X"1000C1000C1000C1000C1000C10006080060840077330C4889CC292588300C00",
INIT_16 => X"44C82082068C0200000008014023EF80020201904189003003000C1000C1000C",
INIT_17 => X"4110441104411044110441104411044110441104411044110441104411044510",
INIT_18 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_19 => X"2FFFFFFFFFFFFFFFFFC110441104411044110441104411044110441104411044",
INIT_1A => X"0924821409005312E8A25E15A69A6BFB0A196A8C5A2932F7C13C15DA08080000",
INIT_1B => X"C46231188C462311892492492492492492492492482082082082082082092482",
INIT_1C => X"00162B158AC562B158AC562B158AC562B158AC562B158AC562B158AC562B1188",
INIT_1D => X"0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"00087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04000",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040200000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"94A7B2B1450000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"6FEBEF5FEC737AFBC6F85FDEB220109E1FEFFFE3FBA7FDFB9BD301DC3FF5F0D2",
INIT_05 => X"FEEDBFDC387F987FEF7C3FAF87FF59F7F5FB7FF59BE1FF980BBBB7FE6D21F3DB",
INIT_06 => X"DFA08957902FFDEE9D7DC9D7DF2B263893479DDFAFDFE15213FFFBE1F1D3A333",
INIT_07 => X"00018010992310605CE10301DE0C1831CB7DF60A244B9BFEE00589DDBCEFEDC1",
INIT_08 => X"FFEFAA001D8EA111DA7FEFF90F21C8C84D9C0D858FC7020828C18FD18346BBF0",
INIT_09 => X"0BFAFFF37DF7B9DF7DCB3FDE89ECC07DF7DF5F985C6BCFFBFA28F99E7EB07F47",
INIT_0A => X"0607307DCFE1D4077B4D0026FFFFBE7D67D7F3BB79CFFB83BF14EC1E7D598058",
INIT_0B => X"FFFCFFC7D7D51D6F5FDCB935D7AFEBD7F5EBFBF7FEBD66DBFCA3F87501AE7B08",
INIT_0C => X"40520201F45EC0010007E01001F45EC0010007E010084BCD7FF1B61B5C33813F",
INIT_0D => X"0001A001F45EC0010007E01001F45EC0010007E01001BD8020500008001F0100",
INIT_0E => X"0200001EC00040B02007EC09A0E00010001DC0004600400F781429C008000077",
INIT_0F => X"81C203404B3BFD0402346235408402C08010003C064000E408010081BD802060",
INIT_10 => X"68B1000E401A08FE0012040000FC002001360403E434588007200D00F88C84C0",
INIT_11 => X"281D00001F01002156040675809145400007B00040091F1190982038406807C8",
INIT_12 => X"903A80008320C0403C34000088601604067D00212000007C400082D81009FC08",
INIT_13 => X"D6BFDFF7BFFED3FBFF6A84383F177FF005FFBFF5FA1040076065F730FC08043A",
INIT_14 => X"CDEBCFF589807B7096CD4CF73AC1FC98884FFF19FFC71FEFED7B251E35768E8E",
INIT_15 => X"78C0D78C0D78C0D78C0D78C0D7A606BC606B8C56F7730ECCDBDF152199F51EDD",
INIT_16 => X"FEFDFDDFE7DD87FEFF7FF796FFFFFDFFD7E681B867D3683A03A40F78C0D78C0D",
INIT_17 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFB",
INIT_18 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_19 => X"6FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_1A => X"4C30C375E2BD54D5D6C565F871C71D44FCF491E166CC853E8695F86EDB5C8864",
INIT_1B => X"26130984C26130984C30C30C30C30C30C30C30C30C30C30C30C30C30C30D34D3",
INIT_1C => X"000130984C26130984C26130984C26130984C26130984C26130984C26130984C",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"1085B0B041000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"6FAB975B6470BAF386C87A9CB00000001FEF9F23E3A7BDE79B5101D23FB5C0C2",
INIT_05 => X"F8EDBFD4347F18778E723F2E47FE59C7F5FB7F759B91FB880BA3B6FE2921CBDB",
INIT_06 => X"DFC00147000FFC128D5CE8D5CC210638A046889CAB57E84217FFE3E181932377",
INIT_07 => X"000141000000042000000288020C18300320620A80231BFE200181092CE7ED80",
INIT_08 => X"FEEF22000C562551D87E8FF90041101042110180004102800008801183468180",
INIT_09 => X"0BE0FC137FF7A0FF75813F1C85244071EFBF17D85C738BE3FA08F9DE36B05B07",
INIT_0A => X"040510768EA0C406630D00226FFE3E2D62D6E21259CFDB039E806C0245188040",
INIT_0B => X"FF48FFCC57550D63564D1D2556ADAB56D5AB6AD7EAB962CBD8A3A83101F47E08",
INIT_0C => X"00130201E44A40010007600005E44A4001000760000843C561E5C55C42B9011F",
INIT_0D => X"00002005E44A40010007600005E44A40010007600004BD8020100008001F0100",
INIT_0E => X"0200001EC00000382006EC0820A00010001DC0000208400D781020C008000077",
INIT_0F => X"81C20040431BC50402146235400400408010003C064000C400018080BD802020",
INIT_10 => X"4821000E400204FE0010040000FC0000003E0403A424108007200102E8888080",
INIT_11 => X"080500001F0100005E040475808101400007B00000015D111010203840081748",
INIT_12 => X"903A8000012040403C34000080201E04047D00202000007C400000F81001FC08",
INIT_13 => X"109E1FE5ADA4C25ADE72041A3F147FF0018DBBB5FA10400360649310FC08003A",
INIT_14 => X"EFABC7054880693016DD4C755AC16C1A884FFE18FFD757E7ED7A211E81C09818",
INIT_15 => X"3440C3440C3440C3440C3440C3C2061A2061AD46FF730E5CCBCD55219AB55F0D",
INIT_16 => X"DE75ED5EC71385FC2512E3565BBBF1BAD6F281BC63F1683803C00E3440C3440C",
INIT_17 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6B",
INIT_18 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_19 => X"7FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_1A => X"0000003C010072F24388521000000140A8100481CA8604368714104A47168874",
INIT_1B => X"8040201008040201000000000000000000000000000000000000000010400000",
INIT_1C => X"00140A05028140A05028140A05028140A05028140A05028140A05028140A0100",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"8C2100804900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"02000100440408002408008002221000204116A280000F000001400000100010",
INIT_05 => X"0004D44400004D4400000000000000000000005C0000000A0000002C20600000",
INIT_06 => X"2000004100000120040A0040A00B009000620294010000400080000888800911",
INIT_07 => X"2488045002489020420110800244891211440804000810002000081040000000",
INIT_08 => X"00B062080542C004CA00000050080202008401842004108AAAA00008912240A1",
INIT_09 => X"2800010000000C0000E400002040500000009202C10020400044000222000204",
INIT_0A => X"02043058C460540329810002D002000400407020800000004000640800088008",
INIT_0B => X"0008000140000401028008330000800040002002480102010082981500062108",
INIT_0C => X"00500000040A40000000A00000040A40000000A0000040060084104110828030",
INIT_0D => X"00012000040A40000000A00000040A40000000A0000000800010000000000000",
INIT_0E => X"00000000000000A00000040020A000000000000006000000080020C000000000",
INIT_0F => X"8000024040152000000020000004004080000000000000240000000000800020",
INIT_10 => X"0821000000120002000004000000000001220000040410800000090000808080",
INIT_11 => X"0805000000000001420000200001014000000000000900101010200000480008",
INIT_12 => X"0000000001204000000000000820020000200000200000000000028800002000",
INIT_13 => X"29400000933050080C0001900020000000408010000000022000D61028000008",
INIT_14 => X"440245400082D022040000400800081022C0000080000206CB0821082B694D4D",
INIT_15 => X"605016050160501605016050160280B0280B0012000843066021001400040024",
INIT_16 => X"0810840861CD33548542A10209D4100E4040A00002002C004001036050160501",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008021",
INIT_18 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_19 => X"0000000000000000000020080200802008020080200802008020080200802008",
INIT_1A => X"41041001A835050788440B58C30C31DF6C110A00246972C0C39989A40A0C22E1",
INIT_1B => X"C06030180C060301810410410410410410410410410410410410410410410410",
INIT_1C => X"00160B0582C160B0582C160B0582C160B0582C160B0582C160B0582C160B0180",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0803B2814D0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"26E1E905CC574828C4F85FC600000016004F77E2F887CDB80BC340DC07D1F000",
INIT_05 => X"FE1DFE4C080F884FE33C078F803F19F011E93ED49BE01F1A03B8972E6D20F049",
INIT_06 => X"64A08857902000DE142D4142D5030010134395D70589415002FFF800F0C38111",
INIT_07 => X"00088400092300601CE00101DE040811D919F402244293FEE00400CCB46BA4C1",
INIT_08 => X"7FA0AA08148A4000887FE0000F20C8C80D080D818FC2000000418FD08142BAD0",
INIT_09 => X"0BFA02E204D2154D28AA3FC60888D03C10415A80402847F8002458926A002E45",
INIT_0A => X"0406305587A1540231410006DFFF80540541619968C76980E914E4163D498010",
INIT_0B => X"FFFC0007C7C0140D0B50A8218102C0816040B1225C1506512C83E85500AC3A08",
INIT_0C => X"40520000141EC0000000A01000141EC0000000A01008480D3EB4A24A0C910037",
INIT_0D => X"0001A000141EC0000000A01000141EC0000000A0100100800050000000000000",
INIT_0E => X"00000000000040B000010401A0E000000000000046000002080429C000000000",
INIT_0F => X"80000340483B590000202000008402C080000000000000240801000100800060",
INIT_10 => X"28B10000001A08020002040000000020013600004414588000000D00108484C0",
INIT_11 => X"281D000000000021560002200011454000000000400902109098200000680088",
INIT_12 => X"000000008320C00000000000086016000220000120000000000082D800082000",
INIT_13 => X"D6ABC032936E43A92F2880B01F37001004B29450580000066021F6303C000408",
INIT_14 => X"45624DB481806A62840800C22800B8900042FF0180000ABFEF89250815568A8A",
INIT_15 => X"68D0068D0068D0068D0068D006A68034680300021410028450530014014002D4",
INIT_16 => X"2C989489418D13FE7F3FFD8BADB7FC4F4164A00806522C0A40A50268D0068D00",
INIT_17 => X"C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C4B1",
INIT_18 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_19 => X"2FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_1A => X"5D75D7FFEFFDF9FAF3E7E3EFFFFFFEBFD6EE7FFDF7FE78FC3CEFFDFFEA0C0060",
INIT_1B => X"EFF7FBFDFEFF7FBFDF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DD75D75D7",
INIT_1C => X"001F7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDF",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"3CF3CF75EFBD75F5FFEFFDFDF7DF7FFFFEFF9FE1F7FFBFEFDFBBFDFFD0000000",
INIT_1B => X"FE7F3F9FCFE7F3F9FCF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"0007F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"1084B030000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"6DA986092050306382C05A1C900000001FAE89016387B2A38B5000D03FA1C0C2",
INIT_05 => X"F8F92B90307F41338E303F0E07FE19C7F1FB7F289B81FB8003A396D20940C3DB",
INIT_06 => X"DF800106000FFC020004C0004C0006288004880800036002137FE3E101030222",
INIT_07 => X"000100000000000000000220000810200220620E00030BFE000181092CE7ED80",
INIT_08 => X"7E4F400000000001107E8FF90001000040100000004102200000801102448100",
INIT_09 => X"23E0FC027DF780DF74013F1C00240071E79F05888C618BA3F800599C10104903",
INIT_0A => X"040100240A808004420400202FFC3E002202021259CFDB039E00080245100000",
INIT_0B => X"FF40FFC407500020004C10060204010200810040801060C04821202001A05A00",
INIT_0C => X"00020201E04000010007400001E0400001000740000803C0616184184031010F",
INIT_0D => X"00000001E04000010007400001E04000010007400000BD0020000008001F0100",
INIT_0E => X"0200001EC00000102006E80800000010001DC0000000400D7010000008000077",
INIT_0F => X"01C200000308C50402144235400000000010003C064000C000010080BD002000",
INIT_10 => X"4000000E400000FC0010000000FC000000140403A020000007200000E8080000",
INIT_11 => X"000000001F01000014040455808000000007B00000001D010000003840000740",
INIT_12 => X"903A8000000000403C34000080001404045D00200000007C400000501001DC08",
INIT_13 => X"001A1FE004048240426200081F147FF0018C1380DA10400140640100D4080032",
INIT_14 => X"812982050800A91012494C31004124080886FE187FC301B124F2001600000000",
INIT_15 => X"1000C1000C1000C1000C1000C18006080060840477330C4889CC012188310E08",
INIT_16 => X"44602002061004A820104809402BE1900222019861D1403803800C1000C1000C",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"2FFFFFFFFFFFFFFFFF8100401004010040100401004010040100401004010040",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000100080",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"88280C4C7B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"00160090920C04800904848262220277E05152B280780D407428E723C01E1400",
INIT_05 => X"0006D46207801E400183C0707800E6000E008057641E00473C40680D32330C00",
INIT_06 => X"203F70C165000225E2C11E2C12A0D0144AC27206582C166504800000B0FC21D5",
INIT_07 => X"920CFC5E6D233B964E7CD99DFB870E1DDDD889C5FBDC440129A0604442180238",
INIT_08 => X"80B036AD23C17544C581000657A0E8E83D86F0E4A7B2D88AAAFD7FE0E1833AC5",
INIT_09 => X"C800016D82082E2081B6C0027ADA398000008A504318404005B70663212C04A0",
INIT_0A => X"4AF4AA414568729139FAD610C00001A2502440888420247041E87681008CE9AF",
INIT_0B => X"00890022B826E250B12346F1244812240912048941621804A150CA1CA45C254D",
INIT_0C => X"B2E0F1F80FA97FE0F0009E0FC40FA97FE0F0009E0FC048211E9C11C31F82E4A0",
INIT_0D => X"C3CB5F040FAB3FE0F0009E0FC40FAB3FE0F0009E0FCC42EFDFBF0AE03080E2AE",
INIT_0E => X"187806013879BA878FE807F65FBF12E0380231F0BD9E3FC08FEBD6F661C0E008",
INIT_0F => X"C83136B248831ACBFC8BBDCAB779BC699F20180309A0F83BE2B87C7C42EFDFBF",
INIT_10 => X"9947184131B59003FFEC07F00003F01FB90BE9F01FC8B38C2098DAE007F323A0",
INIT_11 => X"D065703080E29F1B2BE9F8A27E6E915C0E004C72BEC800FE7464290626D7003F",
INIT_12 => X"6F846DFC0C2352A0024B83F07F198BE9F8A0FFDA2A3C0202B8776A2FA7F023F7",
INIT_13 => X"11800014481A6105810941C5C068000CD4004C0905E52630BB1AE49C2BA7F98D",
INIT_14 => X"7E96656074EA560F0416A24844B01302A26100C4801844069B0C88881A28C141",
INIT_15 => X"E2781EA781E2781EA781E2781C33C0613C0E21020800239450116ED443C041B4",
INIT_16 => X"8112C1241140A056954AB0C280D0002020187007122C3E04E03383E2781EA781",
INIT_17 => X"1204812048120481204812048120481204812048120481204812048120481205",
INIT_18 => X"2048120481204812048120481204812048120481204812048120481204812048",
INIT_19 => X"4000000000000000001204812048120481204812048120481204812048120481",
INIT_1A => X"10410411062084E57CE2641DC71C71574E09B56C74DAB16782171CF13043A85D",
INIT_1B => X"F87C3E1F0F87C3E1F04104104104104104104104104104104104104104104104",
INIT_1C => X"0007C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0",
INIT_1D => X"0000000000000000000000000187C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE500",
INIT_1E => X"BD54BAF7FFD55EF007FD75EFFFAE97555557BD75EF5D00000000000000000000",
INIT_1F => X"FFC0000AA843FE00AAFBE8B45AA803DFEFA28428B455D0017410A28428AAAA2F",
INIT_20 => X"57FFFEBAA2D5401450051401555D7FC0145F7AEBFFFF08002AA10A2AABFEAAA2",
INIT_21 => X"5D7BD755555517FFEFA280021FF082E974AA5D7BFFE000804000BAAAAAAAB455",
INIT_22 => X"A5D2EA8B45005168A10AA8028A10087FD7410557FC21555D51574AAA2FFE8B45",
INIT_23 => X"FFFFAE95410AA80000005D003FEAAFFAEBFE00A2803FEBA002A820AA0800174B",
INIT_24 => X"5EFA2AEA8A10000417410A2FFE8BEFF7FFE8B45FFFBC00005D003FF45557FC01",
INIT_25 => X"000000000000000000000000000000000000000000557DF5500003DFEFFF8417",
INIT_26 => X"12555F524AFE38B780154BAFFF1D54AF0075D75EFEBAE9554540754717F1F800",
INIT_27 => X"B6AB50B6AABDE12BEA0AF010B7D1F8F47E00A2DB45AA8A3AFD7B68E2AB78550E",
INIT_28 => X"A43FE9257F1E816D557095EAAA2D1401D500002A150038038E285D7F78FD7000",
INIT_29 => X"57545A87AAD178A8002D1D21C5E8257D5C7AA854008700249243A412EBFF5542",
INIT_2A => X"02D152A82000E3A5D2150AB8F401471EDBC0B680900AAF52B474385D75C502D1",
INIT_2B => X"D417FD7E9541242FE920AD082E10A28F6A150012A2F02AFFDF40E85F475451D5",
INIT_2C => X"55080550E87B7A405B52AAD152BD00151EAFEDB52E3F1EFFFF485A2DA3D5D24B",
INIT_2D => X"445057F40545850000000000000000000000000000000000000000000005AAF5",
INIT_2E => X"AB55F7AEAABFF5D2A81151FB8635A02FA69574BAF7D5555AF0D79D55FFA2AC97",
INIT_2F => X"34A08D46F6ABE7082AAAAF2FAC77FE00FF16565B2FA9075F4F7B3EBDF50FEAEA",
INIT_30 => X"C95256803CE3AEB038662E5D81406014D5D51F5E08A394003A908B8410E707EF",
INIT_31 => X"C0954AF0151555AF58794040077D774FAE8C798A11A0EAEF75F7AA84001A7052",
INIT_32 => X"245B4E1870108B11020AD4AA05542A0A05051023F9A9D57B63BFBF906CB45FAB",
INIT_33 => X"ABD5F5F0DA6BC9525688C1A2A0C06E9FEE5555BE48AB2A2AE0A0F20C43EAC562",
INIT_34 => X"0FF8000000FF80F55E25C00A0BA7FBED407A97F6F35F498B96BEB12DAAB77558",
INIT_35 => X"00FF8000000FF8000000FF8000000FF8000000FF8000000FF8000000FF800000",
INIT_36 => X"000000000000000000000000000000FF8000000FF8000000FF8000000FF80000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000800000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"CA1800080848B0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000010822C00803804000001999EF9C00040B0002000001000640200001018",
INIT_05 => X"0000400244000000014200004000000004000000001000032000200002100800",
INIT_06 => X"202800208500000080412804100CB08000302220080408010000000404100844",
INIT_07 => X"25FC4C5AF6FEF002230018010860C1833C460044204C000008A0041000080008",
INIT_08 => X"0010008D22C0F55000010000524481890BC000263000188AAAA10F8C1830562B",
INIT_09 => X"041001B102002E20013600022D8819000000A000110A4000002C204000240420",
INIT_0A => X"0BE0B002605C1C1108484400C000002040040820000020104100028800002801",
INIT_0B => X"000000081001004010810510040802040102008100200800A1100707040101E2",
INIT_0C => X"10F18058000003C0F000A000C4000003C0F000A000C0000012187087010AE4B0",
INIT_0D => X"00012704000003C0F000A000C4000003C0F000A000CC4200002F08E030800000",
INIT_0E => X"1878060000000AAC00680000001F10E038000000078808C00000023461C0E000",
INIT_0F => X"4800025200040A00D000000202090C281F201803000000240218C0044200001E",
INIT_10 => X"904618400012900001EC03F000000000392100B00048230C200009A000130320",
INIT_11 => X"806070308000000961002880204A901C0E00000002C9000260640900004D0000",
INIT_12 => X"0904285C0C0312A002000000083881002880025A0A3C020000002A8400B00007",
INIT_13 => X"08400004080030008010468220A00008D0000801046004308A18500002012800",
INIT_14 => X"2200000840280206089000004090110200000000001454000200828008081110",
INIT_15 => X"A4191A4191AC191AC191A4191A00C8560C8D2910000060901010401E13405111",
INIT_16 => X"8000410410028000100800140000002004103224002006406401918C191AC191",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"0000000000000000000200802008020080200802008020080200802008020080",
INIT_1A => X"1451455901218D2C4CA2900C9249258306BABEFC54A081701C397452B4008A04",
INIT_1B => X"BADD6EB75BADD6EB755555555555555555555555555555555555555545145145",
INIT_1C => X"0005D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2EB75",
INIT_1D => X"0000000000000000000000000607FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF600",
INIT_1E => X"E80010AAAABFFFFFF803FE10F7D17FEBA55556AAAAAA80000000000000000000",
INIT_1F => X"2EBFEBAFFD555400557BD54BA5D7FFDF45A2FBD75EFA2AE97555F7FBFFF45FFA",
INIT_20 => X"A802ABEFA2D568A005D5157400AA8028AAAF7FBD54AA002A955555D7FE8ABA08",
INIT_21 => X"FFFFFDF55AAFBC0010555540010550417555AA8028BEFAAAE97555082A80000A",
INIT_22 => X"A557BD7410550428ABA5D5168ABA552EBDFEF5D7FEAA00AAAABFEAA007BC0145",
INIT_23 => X"FFFFFFEAB55557FFFEBAAAD568B45A2D5575555D7FC2155F7AEA8BEFAAAA954B",
INIT_24 => X"4AA5D7BD74000804154BA082ABFF55FFD57DF45F7D568ABAF7AABFFFF082ABFF",
INIT_25 => X"0000000000000000000000000000000000000000002EBFFEFA280021FF082E97",
INIT_26 => X"95545E175EFF57BF8FC2000BEA4BAE97F78A3FE28E3D17DEAA485FE8E02B5000",
INIT_27 => X"FD55455571E8A2A087BF8EAAEB8E0016D5D75D54BA5D7BFFF7DA2FFD55EFAAA4",
INIT_28 => X"AA07157428145A00AA8A2FBD7B6DF6AA28550E10405F7A4AFE38EAA0924921C2",
INIT_29 => X"6AAB8E971471C7010B7D168F47400A07A28415A001684104155C5B6DF6DBEFBF",
INIT_2A => X"5FD4BFBD7B6A0BF492415FC20105D24AAABF1FFBC7010FF8A38FEF557FEAB78B",
INIT_2B => X"FE38017EBA4A8EB8F6FFD5FE8B7D557495EAAA2D16D1FDBED56A55557A43DE38",
INIT_2C => X"C7AA854008700249243A417FFF41542F5D717FE2AAAA56DEBD17FE3DF7FB7FEB",
INIT_2D => X"FBA007DFCA127B8000000000000000000000000000000000000000000002A3D5",
INIT_2E => X"FFEFAAFBD55FFAA8416545A6FB60F47AF2A00010F78028B15F7823FEAAA2D57D",
INIT_2F => X"21A022A38C20B2552E975F758516AAAA0869AAAB8A7C19C55550E8574BA557BF",
INIT_30 => X"895755FFEFBCEE5FBAACB10085EE5DE10A2AEBFF55F7BAAA8565DBAC1112FFAC",
INIT_31 => X"02EABEA097BEAAFAF2863FA00DD574201E7AD1FFF5575841DE08007FC2048002",
INIT_32 => X"AF9554FF57EFBFA18D4FBFFF40FF809D4000D7FC00FC5D062BBA05ED5034472A",
INIT_33 => X"FED17DFBFF6963FCAAA2283CF14050062B0A2F7AE8B5D5D51F5E18ABD5EAFFF2",
INIT_34 => X"0000000000002CB75F7AA84001A7052C95256807DC31AA8114DE55F5BED201FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000800000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E44660018259B2843913100062C98004802322D3E030235201006009B2812",
INIT_01 => X"0005A18A0849204D1CA024A542500368404000720885800802000106E4D10204",
INIT_02 => X"5C010802020408040C600850AA055254090541A111240A104A0000000908B510",
INIT_03 => X"182202210800004401060A0010041028021560A0218808002440840008C80550",
INIT_04 => X"21030A008814500120A06B0870201010258261E141A2326511024182142494D2",
INIT_05 => X"48484098142953388552102442884882B58A09291290A1120A81A3C200418DCA",
INIT_06 => X"22208802800554529001C9003A2800203120000104810100002A614008102244",
INIT_07 => X"0008040000221040408100890C0000011804480420420154000088096A0EA8C0",
INIT_08 => X"B846C0081190C105424705510A08828A0B190C0428040080A0A10F8000009200",
INIT_09 => X"20B0573165541CD54822160A89E89020AA8A80CA9D39CE215264B15818004442",
INIT_0A => X"0402100C088104010AC80005C568147007031012D40D71824114081538000048",
INIT_0B => X"550055481205100C000134128304408020C11020040244D00001306100A24600",
INIT_0C => X"00500000B01480010000A00001501480010000A0000801487334E34C1A980001",
INIT_0D => X"00012001501480010000A00000B01480010000A0000138000040000800000000",
INIT_0E => X"02000000000000A00003600180400010000000000608000A5004090008000000",
INIT_0F => X"000002400008C4000220420040800280001000000000002400000001A1000040",
INIT_10 => X"2090000000120C94000200000000000001380001C01048000000090298040440",
INIT_11 => X"2018000000000001580002508010440000000000000953008088000000481380",
INIT_12 => X"10180000820080000000000008201800024C000100000000000002E000095000",
INIT_13 => X"09130A82000C90A0000081A004342AB001720040000000000001502050000422",
INIT_14 => X"094882958000934200904407600090822085E0100D52498002B1041092001514",
INIT_15 => X"3C1011C1013C1011C10134101140801A0808AD4451394CD0391A541593C04B59",
INIT_16 => X"022810800000A0289A6D084D4021208106142034406144004041011410114101",
INIT_17 => X"4010040104411044110441100401004010040104411044110441100401004010",
INIT_18 => X"0102401024010241106411064110640102401024010441104411044110040100",
INIT_19 => X"2F81F81F83F03F03F04110641106411064010240102401024110641106411064",
INIT_1A => X"0820823047486021658010816596597700138D70C030B542923650C7D0002281",
INIT_1B => X"944A25128944A251282082082082082082082082082082082082082082082082",
INIT_1C => X"F804A25128944A25128944A25128944A25128944A25128944A25128944A25128",
INIT_1D => X"0000000000000000000000000787C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF871",
INIT_1E => X"5420AAAA843DFFFAAD1554005D7FD74AA0004001550000000000000000000000",
INIT_1F => X"2EBFF45AAAAA8A10A2AE80010A2AA975FF5D003FE10F7D17FEBAF7D5420AA085",
INIT_20 => X"D7FFFF45A2AA975EFA2FFD7555FFFBFFF45AAFBC20AAF7D1575EF55517DF555D",
INIT_21 => X"AAAE95555552E974105D517DF55AAAAAABEFAAD1575EFAAAE974AA5D51554BA5",
INIT_22 => X"F552E82010F7AABFE10FFD542145FFD5554AA555555555557FE8ABA082EBFFFF",
INIT_23 => X"EFF7FBC0010AA802ABEFAAD540000FFD540000AA802AABAF7FFC2010AAAE821E",
INIT_24 => X"555AA8028BEFAAAE821550851420AA002E800AA08042AB45007FC00BAFFD168B",
INIT_25 => X"0000000000000000000000000000000000000000002E80010555540010550417",
INIT_26 => X"7DEAAE95F40002157F470AABE803AE97A2DF55400557FD54AA1D04001C515000",
INIT_27 => X"E105EF55517DFC5552ABDF45B6AEAFFD5F7A482000BEAE905C755003FE28E3D1",
INIT_28 => X"A4070BA5FD0154BA5D7BFAF7DA2AE955EFAAA495545E3F5EFF57F7FE80082FFD",
INIT_29 => X"571E8AAF082AB8EAAEB8E0016D5D2A924105D5B7FF7DB6AAAABC7BEDB505EFBE",
INIT_2A => X"E80495038AAAEAF1D7410E80000FF8438E00B6DF68FEF4871D24BA495B5556D5",
INIT_2B => X"80071ED1EFEAF1EFFFDEAD1C5010AA8E2FBD7B6DF47A00EBDB50000A380AAE28",
INIT_2C => X"28415A001684104155C5B68E2DBEFBFFBC703AE2DF42AAA002A851C214003FF6",
INIT_2D => X"4AA550002155510000000000000000000000000000000000000000000002087A",
INIT_2E => X"215555003FEAAAAD57DEBAA2FDDC01051FBD74BAF7802AB05AAFBD5400557BD5",
INIT_2F => X"60F47AF7FC20B2F7FBC015D58517FF555D2ABDF55F782BEB47AFAD00010F7AA8",
INIT_30 => X"22A955FFFFC20FFF3AE544108410174BA557BEABEFAAEBD55FFAA1456547A2D3",
INIT_31 => X"D4420BA547FD75FF58516AAAA0828AAAB4A78016545540400010557BFDFFFF78",
INIT_32 => X"FFBD550AAFACAAA122AA8954BAA2AE9D545002A800A8FF862BA00F2F9E8F0050",
INIT_33 => X"002E954505C417FFFF08555555BAAD335B57AB5155400A2AEBFF45FFFB404007",
INIT_34 => X"000000000000061DE08007FC2048002895755FFAEBCFE57BBA57002DF3C4AAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000001000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C00A20020000108430020001600B815602110494074133520400E02B92206",
INIT_01 => X"014C9BC048800168240442C99E004B61404040028804A0080A000516A0990A08",
INIT_02 => X"4809A900031800444440589866E331352180D468B8000E600C0081110B802CD0",
INIT_03 => X"DA16C0200C0001423583480408D60520320066810A80881068A808029C856330",
INIT_04 => X"2088681DA82740EC92307364B37569100A84E1E11C251210990040420E005A48",
INIT_05 => X"2D284A102414411A314A0A02C18C01B9854368280A506902018C2442484038D1",
INIT_06 => X"23600016801CCCAA9061C9061C0D0080001005210C8761001166CCC40C110826",
INIT_07 => X"0178045800B6540063000889082040A13A0716042440833280038C89904E6400",
INIT_08 => X"D20A480810804451421D1CC8024481994B5500061000088000A10F840854973A",
INIT_09 => X"2079CCB035E03CCC5D2A35620988100A698761C0953B6E84C82C404018304D42",
INIT_0A => X"070070202A90340440C80004CCE4CC1042061913208CE8024380880820010040",
INIT_0B => X"3302CCC01300104018900402870C4287214210E114200410EC20242D01015E84",
INIT_0C => X"4801000180148000000800100040148000000800100401C33249049051218073",
INIT_0D => X"04008001001480000008001000E014800000080010001C000040000000000000",
INIT_0E => X"0000000000004408000068018040000000000001400800091004090000000000",
INIT_0F => X"00004100812644000004400140800280000000000002000008008000B0000040",
INIT_10 => X"20900000020800CC0002000000000020400800030010480000010400C8040440",
INIT_11 => X"2018000000000060080004418010440000000000410015008088000008200540",
INIT_12 => X"80188000820080000000000100400800041C0001000000000000902000014C00",
INIT_13 => X"284B264208448260E27285A23224E660084208410000004444000E0000000020",
INIT_14 => X"0840024D810283021280400720C0348002854C001CC3158026A2040028090441",
INIT_15 => X"80901A0901A09018090188901A248054480C0C0041116DD0115E011599641E59",
INIT_16 => X"C6C8408514028028D06C0C5D20030BA1010021B000020402400501A090180901",
INIT_17 => X"4290C4290843908439084390843908439084390C4290C4290C4290C4290C4690",
INIT_18 => X"290C4210E4290C4310A439084310A439084310A4390C4290C4290C4290C4290C",
INIT_19 => X"5D54AAB556AA9556AAC310A439084310A439084310A439084210E4290C4210E4",
INIT_1A => X"0820825103A1600054C0F4012492490300C78C706428A1411133586294020A90",
INIT_1B => X"D4EA753A9D4EA753A92492492492492492492492492492492492492482082082",
INIT_1C => X"8086A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A353A9",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE024",
INIT_1E => X"5421EFAAFFD54AAF7D168B45AAAABDF5500002AA100000000000000000000000",
INIT_1F => X"043DF45FFD168AAA0855420AAAA843DFFFAAD1554005D7FD74AAA28400155005",
INIT_20 => X"2AA955FF5D003FE10F7803FEBAFFD5420AA080400155AAD5554AAF7802AB4500",
INIT_21 => X"AA8028B45A2AE82155A2FBFFEBA0800021550855555FFAA84001FFAAAE80010A",
INIT_22 => X"0085168ABAFFFBD54BAAAAE97400A2FBC20AAA284175EF55517DF555D2EBFE00",
INIT_23 => X"55AAAA954AA5D7FFFF45AAAA975EF007BD7555FFFBFDF55AAFBD55EF5D2EBFE1",
INIT_24 => X"BEFAAD1575EFAAAE974AA5D00175555D0015410F7AAAAAAA55043DE00FFFFD55",
INIT_25 => X"00000000000000000000000000000000000000000004174105D517DF55AAAAAA",
INIT_26 => X"D54AABC04001C51551471D7AAF1D05D2EBD56DB7DBEAEBFF551C042AA101D000",
INIT_27 => X"B50492EB842FB5508043FF55EBD56ABD75D5B470AABE8A3AFD7A2DF55400557F",
INIT_28 => X"8E82557FD2082000BEAE905C755003FE28E3D17DEAAEBDF40002550F47155AAD",
INIT_29 => X"5517DF40552ABDF45B6AEAFFD5F7A48017DAAFFFAE821C0A0717D1C5B575FFB6",
INIT_2A => X"F7D5C55D7492E90E3808756DA92EBFFD74BAE3AE85480FFFFC00AABE8E105C75",
INIT_2B => X"241043AE10EAF5C5547FF80954AA5D7FFAF7DA2AE905EF0075D5545E3F5EFF57",
INIT_2C => X"105D5B7FF7DB6AAAABC7BEDB505EFBEF5C7092FF801756D490A10438EBA4B8E9",
INIT_2D => X"F555D0028A00510000000000000000000000000000000000000000000000E124",
INIT_2E => X"8B45AAFBD54005D7BD54AAF78002155515157555AAD142040A2D57FFFFFFAEBF",
INIT_2F => X"DC01051AE955F7AAFBC0000AF843FF5500003FF55AAFD6AB455157D74BAF7AAA",
INIT_30 => X"E955FF557BD74EFFBACD41577B8400010F7AA8215555003FEAAAAC53DEB8A2FD",
INIT_31 => X"FEC20BAF7AA8015558517FF555D2ABDF51F782BCB47ABAE801FFAAFBEAA105D2",
INIT_32 => X"8554214FA2D3EAF57AFFDD7555082AA0AAA00557FEA8A2FDD64BAAF8282012AF",
INIT_33 => X"082A820AAAB842AA00000028AB0AAFF48547AE04174BA557BEABEFA2AA951FF8",
INIT_34 => X"0000000000002A80010557BFDFFFF7822A955FFFFC21FFF3BE40412DE02955FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000800000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303000048B3532C82D04A16002",
INIT_01 => X"210399800808004C1C20650E1E104368403008418984014902030006A8910200",
INIT_02 => X"480108A200000000444148E41E80F00A4104311868200200080000000988A390",
INIT_03 => X"0CA08220080000D004260A0240109028270012603000000030808C4208C000F0",
INIT_04 => X"4403A609A055306BC2C0735810CEE5100A0A48E16B8370E3808241D03845D002",
INIT_05 => X"ECE8698800791403AD3038AE079059A790E245A19A41E4120BAB86C00001D312",
INIT_06 => X"23208806000C3D220023C0021A21008891048C00040341121661E3C10000A064",
INIT_07 => X"0008045000220440000000090800102118400204A04100F040018019004B8001",
INIT_08 => X"0E11400810906441123323C0424190880B0108002000000880810F9002041200",
INIT_09 => X"22003C2309671584786E0F5A88889031EF9F05D884794FA03A24781810106D02",
INIT_0A => X"0409400E4282A00142400004DC3C82400702003200872003FB14080828400010",
INIT_0B => X"F050C3C00095000C008135040002010100800040001400C00401208800F01A14",
INIT_0C => X"08000002E0100000000800000220100000000800000001C87261C51C42390240",
INIT_0D => X"0400000280100000000800000360100000000800000035100040000000000000",
INIT_0E => X"00000000000004000000D8008000000000000001000000155000080000000000",
INIT_0F => X"000040000120EC00004002214000008000000000000200000000000094100040",
INIT_10 => X"001000000200050C000200000000000040080005800008000001000168000040",
INIT_11 => X"000800000000004008000448000040000000000001003C000008000008000D00",
INIT_12 => X"800800000000800000000001000008000017000100000000000010200002C800",
INIT_13 => X"150F5E0400101000227200800E271E00288400800208004C04C0080000000052",
INIT_14 => X"818082450000920280C544310041B408880EC51060461589225100063E9012D6",
INIT_15 => X"1410C3410C1410C1410C3410C100869A08618C00772201D899BA003591510A59",
INIT_16 => X"44E0110004480020986D4815044369A00006203041C3443043010C5410C3410C",
INIT_17 => X"0080001002008040100200800000060180000006008000100600804000020180",
INIT_18 => X"0000010060080201800000040100201802008040100201804000020180001006",
INIT_19 => X"64B261934D964C32698080401000000060080601800000040000201806008000",
INIT_1A => X"1451457A604C8D0C28A280CD145144C1863807E0500014385DAF345041488280",
INIT_1B => X"1A8D46A351A8D46A355555555555555555555555555555555555555545145145",
INIT_1C => X"1F60D068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D06A35",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE077",
INIT_1E => X"02ABFF087FFDF5508003FEBA087FD54BAAA84154005500000000000000000000",
INIT_1F => X"2EBFF5500003DF455555421EFAAFFD54AAF7D168B45AAAABDF55A2802AA10000",
INIT_20 => X"A843DFFFAAD1554005D7FD74AAAA840015500002AABA082E954005500021FF5D",
INIT_21 => X"FFD168BEF080028BFF0855555455500174BAA2AABDE0055517FF555555420AAA",
INIT_22 => X"0085168ABA0055574BA5555554BA5D0400155AAD1554AAF7802AB4500043DF45",
INIT_23 => X"AA5D0400010A2AA955FF55003FE10F7803FEBAFFD5420BA085168A00007BFDE1",
INIT_24 => X"1550855555FFAA84001FFAAFBEAB45002A97545F7D1555EF55043DF5555517DE",
INIT_25 => X"0000000000000000000000000000000000000000002A82155A2FBFFEBA080002",
INIT_26 => X"BFF55BC042AA101D0A28BC7007FFDF45080A3AEAA007BD2482BE84124285C000",
INIT_27 => X"4974004100021FF492AB8F7D1C0438E381451471D7AAFBD0492EBD56DB7DBEAE",
INIT_28 => X"557AFED1C5F470AABE8A3AFD7A2DF55400557FD54AABE84001C5550A28ABA142",
INIT_29 => X"B842FB5508043FF55EBD56ABD75D0428BEF005557545490012482B6A0BAE2849",
INIT_2A => X"557F6DA101475FDE10145F68A921C55504924955524AA140E0717DAADB50492E",
INIT_2B => X"F5D043AF6D405F78E3A1C2002000BEAA905C755003FE28E3803DEAAEBDF40002",
INIT_2C => X"7DAAFFFAE821C0A0717D1C5B575FFB6DF425575D7BEFB55002097555FFD5401E",
INIT_2D => X"010F784000AA5900000000000000000000000000000000000000000000020801",
INIT_2E => X"2000A2D57FFFFF7AEBFF55FF8028A00512EAAB45007FFFF55082EA8AAA087FC2",
INIT_2F => X"02155512AAAA085D04174100800021FF002EA8BEF5D0428ABA595557555AAFBC",
INIT_30 => X"402000FF802ABAA04552ABFF597FD74BAF7AAA8B45AAFBD54005D7BD54AAF780",
INIT_31 => X"2F955FFAAFBC0000AF843FF5500003FF55AAFD6AB4551002ABEF005555555000",
INIT_32 => X"A843DEB0A2FD5600051537DE005D557DE005D7BE8AA85555400100879560AA59",
INIT_33 => X"000417545FFD5421FF5D0428BEF0079FCABA598400010F7AA8215555003FEAAA",
INIT_34 => X"00000000000004001FFAAFBEAA105D2E955FF557BD75EFFBBCD415521FBFDF45",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000001000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DB0A0791B1B41694368283C81F9996A091A32152007AB37B20E07C0C1E002",
INIT_01 => X"881FBC449030884C446A00000034824841280A00084000C8C212812EEA953231",
INIT_02 => X"C809AD5CB118E640A4F408FC011FF0002080000082CCC66609DB7DDDCB1F2036",
INIT_03 => X"4A100E4D3E4C90D290831C824A4204720B20048A88800000B8E0F91028C5500E",
INIT_04 => X"00144884922644001914830051110A71E03040F0105B001C662AE22DC08A3408",
INIT_05 => X"120340220B88820041CDC451B860A6506BEBD08265AE105714505F0152122449",
INIT_06 => X"207F7890752C037372A1D72A398CD084C890EA2950A37E270660182C0D2C8080",
INIT_07 => X"9378355E64B66F96231CC81D2DAB468D38C601C5FFF54FF1C9A46490261C4B39",
INIT_08 => X"7F105CAD1089654115814FC60284A1A93B46F4621030C800001D7FA56891162E",
INIT_09 => X"E00A003C832D25328526C082DF9AB88C104024C09639441807B78661090C24A1",
INIT_0A => X"4FD32A2E2A9992944AF2D611C3FC01B2152109204C28B67061EC928920C569E7",
INIT_0B => X"F0313FE92C22F21CA0B363C0A242502028901408154218144D712664A5F15AC1",
INIT_0C => X"B2F0F1E01BE53FE1F000BE0FC41BE53FE1F000BE0FC80020130841840308653F",
INIT_0D => X"C3CB7F041BE1BFE1F000BE0FC41BE1BFE1F000BE0FCD806FFFAF0AE83080E2AE",
INIT_0E => X"1A7806013879BAA78FC103FF5F1F12F0380231F0BF9E3F02A7FFD63669C0E008",
INIT_0F => X"483136F200A822CBACAB9DDEB7F9BC291F30180309A0F83FE2B87C7D006FFF9F",
INIT_10 => X"D1C6184131B7980DFFFC03F00003F01FB931E9C1DBF8A30C2098DBE2FF7F2320",
INIT_11 => X"F060703080E29F1B71E9F6427EFE901C0E004C72BEC95FEF64E4090626DF15B7",
INIT_12 => X"EFAC6DFC8C0312A0024B83F07F3991E9F21DFFFA0A3C0202B8776AC7A7C9CBFF",
INIT_13 => X"88F4C1C64044A264601144C5F1787E1C812A510885C56620590350ACD3A7D5B7",
INIT_14 => X"9054204DF56A974F92C3E20F24301300082C38C4184F10281204888298284616",
INIT_15 => X"A238CE238C8238CE238CA238CC11C6411C670C10EB4124C2B3923BF5C9710C59",
INIT_16 => X"276A11A03444922898494C5504008401230E71B3100C1634E3138C8238CC238C",
INIT_17 => X"5094650142511405194450942511425114450944519425114250144519405194",
INIT_18 => X"0944509465114251146501465014051944509445094051942501465014051940",
INIT_19 => X"2124B2DA6924965B4D5094450940519425014650142511425014450944519405",
INIT_1A => X"7DF7DF6FEFFCFDFD796ED1DCF3CF3DF6CE7F7B9DB7FF3A7E1FBC6DB7E8418A88",
INIT_1B => X"EEF77BBDDEEF77BBDDF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF",
INIT_1C => X"024F77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDD",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE056",
INIT_1E => X"5574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF80000000000000000000",
INIT_1F => X"D16AABAF7AAA8BFFAA802ABFF087FFDF5508003FEBA087FD54BA080415400555",
INIT_20 => X"AFFD54AAF7D168B45AAAABDF55AA802AA1000003FEBA00002AABA5D2EBFEBAAA",
INIT_21 => X"00003DE005555575EFA2D142145A2FFE8B45FF80001555D2E955FFFFD5421EFA",
INIT_22 => X"F5D7FC00BA5D5568AAAF7AAAAAAAAA802AABA082E954005500021FF5D2EBFF55",
INIT_23 => X"BAFFD5420AAAA843DFFFAAD1554005D7FD74AAAA840014500517FFEF007BEABF",
INIT_24 => X"4BAA2AABDE0055517FF555504154BAA2FBEAA105D2E97410FFD16AAAA5D2ABDE",
INIT_25 => X"0000000000000000000000000000000000000000000028BFF085555545550017",
INIT_26 => X"D24821E84124285C51574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7800",
INIT_27 => X"428A925D2AB8EBABEDB6AA92F7AAA8BC7B68A28BC70075FDF45080A3AEAA007B",
INIT_28 => X"2A925FFFFD1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA105D0A38EBA1C0",
INIT_29 => X"100021FF492AB8F7D1C0438E38145B575EFA2DB45145B6F5EFB6DF78E0514555",
INIT_2A => X"55517DFC70875EABC7557FC20AA415F68AAAF7AAAAA82BE8A28A921424974004",
INIT_2B => X"0FFDB6FABA542ABAE2AF7DF470AABE8A3AFD7A2DF55400557FD54AABE84001C5",
INIT_2C => X"EF005557545490012482B6A0BAE2849043AFED1C0E10492B6FFEFA105D2A9541",
INIT_2D => X"E005D2AAABEFFB8000000000000000000000000000000000000000000000428B",
INIT_2E => X"FF55082EA8AAA087FC20105504000AA5955554BAFFAEBDE10F7FBFDEBA007BFD",
INIT_2F => X"28A00512AA8AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3AAAAB4500557",
INIT_30 => X"57FFEFFFAA97545552A821EFFBD557555AAFBC2000A2D57FFFFF7AEBFF55FF80",
INIT_31 => X"AAAAA005D04174100800021FF002EA8BEF5D0428ABA597FD55FFA2FFD5555FFD",
INIT_32 => X"D7BD54AAF7800015551517DF45005168B55557FC0012087FEAABAF7AAAAA10F3",
INIT_33 => X"FFFFFFE005D2A95410F7FFFFEBA5D2EA8ABAFBFFD74BAF7AAA8B45AAFBD54005",
INIT_34 => X"000000000000002ABEF005555555000402000FF802AAAA04452ABFF592E80010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000006000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0061A01002840002C030028180004003220200403302301C0381A0082",
INIT_01 => X"A74041C838394848188160000C42426041000000090800090210000008510200",
INIT_02 => X"080108200C1000004465580000C0080100000000010432400800800009882050",
INIT_03 => X"080200010C234040842248600210812183806584488000103080014E88C10000",
INIT_04 => X"0040584288A6C210003120000000001002A0E8A910A072101000400A00203040",
INIT_05 => X"04096A019400C118414A00014000002014100128005004020010A0C044C02800",
INIT_06 => X"20200A301223FC029931E9931900002224240249A6D3E808D51FE00909108222",
INIT_07 => X"0008040000220001820000010C0810211A440014A040200E8240089000080002",
INIT_08 => X"0040081A08944010007FA038020080880B0104182000000000090F8102041320",
INIT_09 => X"17E2FD200240B4A409223F020888100808200450001A401BF82C21185C81744A",
INIT_0A => X"0602A0244285180542402180D001BE1907939120000020044184890800011000",
INIT_0B => X"0F0400091081190E4490A502D2A36951B428DB14A688051A5E21214601A01A22",
INIT_0C => X"455D0018101480000000A01034101480000000A01033A0081300000000001880",
INIT_0D => X"0001A0F4101480000000A01034101480000000A0103142000040000000000000",
INIT_0E => X"00000000000041E8002900018040000000000000466800C20004090000000000",
INIT_0F => X"0000034D242C2000502000000080028000000000000000240946800142000040",
INIT_10 => X"20900000001A60F0000200000000002007F000322010480000000D1A00040440",
INIT_11 => X"2018000000000025D00008958010440000000000403F4000808800000068D240",
INIT_12 => X"101280008200800000000000086670000CC0000100000000000087C000301400",
INIT_13 => X"C8B5800720849A72700094A2202301F05103202420000810C219500150002800",
INIT_14 => X"81088A454110030212C140813204D0A0888C000118471DE126805432A62A1586",
INIT_15 => X"4096C4096C2096C2096C6096C444B6004B600C446B0104D09190013589701C11",
INIT_16 => X"108D19D1804A8000904C421852240821978221B0044245B25B456C0096C0096C",
INIT_17 => X"69DA368DA1695A568DA3685A1695A768DA3685A569DA768DA1685A569DA76C5A",
INIT_18 => X"85A569DA1685A369DA5695A368DA169DA7695A168DA3695A5695A368DA3695A5",
INIT_19 => X"7638C31C71C718638E685A569DA7685A368DA5695A768DA1685A7695A168DA36",
INIT_1A => X"1C71C73B676CEDED7DE2F4DDF7DF7DF7CE7F8FF0F4FA957FCF9F7CF7F40A0010",
INIT_1B => X"FE7F3F9FCFE7F3F9FC71C71C71C71C71C71C71C71C71C71C71C71C71C71C71C7",
INIT_1C => X"2BE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"0000000000000000000000000607C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF019",
INIT_1E => X"43DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFF80000000000000000000",
INIT_1F => X"D17DEBA0855421455555574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFF8",
INIT_20 => X"87FFDF5508003FEBA087FD54BA000415400550428AAAAA84021FF007BD54BAAA",
INIT_21 => X"F7AAA8BFFAAD1554BA002A95555A28417400AAFBE8ABAF7FFD54AAAA802ABFF0",
INIT_22 => X"0FFFBD5545080417555A2D17FE1000003FEBA00002AABA5D2EBFEBAAAD16AABA",
INIT_23 => X"FFFFD5421EFAAFFD54AAF7D168B45AAAABDF55AA802AA100000001EF087FEAA0",
INIT_24 => X"B45FF80001555D2E955FFFF843DEAAA2803DFEF0855401FF082EA8B555D7FC21",
INIT_25 => X"00000000000000000000000000000000000000000055575EFA2D142145A2FFE8",
INIT_26 => X"6FA92552AB8FEFF78E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FF800",
INIT_27 => X"E001EF147BD2482BED57AE921451421555551574BAB68A2DA00FFFFFFE38085F",
INIT_28 => X"FFD24BAB68A28BC70075FDF45080A3AEAA007BD24821C04124281C0E2DA82BE8",
INIT_29 => X"D2AB8EBABEDB6AA92F7AAA8BC7B6D5524AA14209557DA28E15400BEF1EFA92FF",
INIT_2A => X"5D0E071FF0071EDA38F7F1D5555000417545B6D178E281C0A38EBA1C0428A925",
INIT_2B => X"70824A8B555C7FC2147F7D1471D7AAFBD0492EBD56DB7DBEAEBFF55BE842AA10",
INIT_2C => X"EFA2DB45145B6F5EFB6DF78E05145552A925FFFF8E3DE82BE8E38FFF0851401C",
INIT_2D => X"000557FE8A00F38000000000000000000000000000000000000000000005B575",
INIT_2E => X"DE10F7FBFDEBA007BFDE005D2AAABEFFBAABDFEFAAFBC00BA007BC0000FFD542",
INIT_2F => X"000AA592ABFE00F7AA821FF557FC0010F7D168A105D55421455155554BAFFAEB",
INIT_30 => X"E95410F7D57DE00FFFBC00AAFBAAAAB4500557FF55082EA8AAA087FC20105504",
INIT_31 => X"2AA8AAA5D0028A005D2AA8ABAF7FBE8A00FFAEAAB45F3D5400BA5504155EFAAA",
INIT_32 => X"7AEBFF55FF8028A00512E975FF08557FEAAF7D157545080417545F7D56AAAA59",
INIT_33 => X"F7AAAABEF005542155000028B555D7FC2145F3D557555AAFBC2000A2D57FFFFF",
INIT_34 => X"0000000000007FD55FFA2FFD5555FFD57FFEFFFAA97545552A821EFFBAABDE00",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000004800000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C02450418800002300500030B313300C418992006",
INIT_01 => X"A34009C0383848481C00E0000E01426040000000080000080200010000510204",
INIT_02 => X"4801082048100000446558000080000041000000000622400800000009000010",
INIT_03 => X"080001038CA14840842248400210812102000400088000003080014688800000",
INIT_04 => X"000040048106000040120000000000100220C8A5108032140004500800603000",
INIT_05 => X"04096A009000410041480081000000201000012800400022801080C0C0C82000",
INIT_06 => X"232086381A8001220021E0021803002224240248040360889100100909000222",
INIT_07 => X"0008055000220409020000090C0810211A04001420602000D2500810000C4903",
INIT_08 => X"8040491A809041100001400042409098090006102000000000010F8102041320",
INIT_09 => X"340C013102002420012200820D89140800004010900A4010002C8118D0024412",
INIT_0A => X"A221A5000800914000400888C00100200B0310200008B2066313894800631400",
INIT_0B => X"0010000800010004088105020100008000400120800000200404002450004000",
INIT_0C => X"4409081C1000000000F001F02C1000000000F001F021141A12000000000010B0",
INIT_0D => X"383480CC1000000000F001F02C1000000000F001F023420000000004C3201C51",
INIT_0E => X"00019860078641084039000000000002C0E00E0E404900E200000000000B0380",
INIT_0F => X"120C8908146000105120000000000004004160C0301D07001D04820342000000",
INIT_10 => X"000021908C4842FC000000030F000FE00600103BA0000010C8462414E8000006",
INIT_11 => X"000004C3201C60A400100DD5800000013098038D40309D000000C2419120A740",
INIT_12 => X"901A800030040902C0807C0E00C440100DDD000000411C81078884004035DC00",
INIT_13 => X"140A000410401400201020820022000250400040002211148019064200402A32",
INIT_14 => X"01889A4543148282A01415B04009904A80890033679459A926801054001C0050",
INIT_15 => X"159201592055920559205592070C901AC901A100804000801210541403C05130",
INIT_16 => X"2460010004428008904C085D44200D8001112804CDE1C483480D201592015920",
INIT_17 => X"0080200806008020000000004000020080200802000000000000000008020480",
INIT_18 => X"1000008020080000000000020080200000000000080600802008000000400000",
INIT_19 => X"5841040002082080000180200000000020180200800000000100200802000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000005428A94",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"E480000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE031",
INIT_1E => X"BC00AAF7D5575455D557DFEF002AAAB55002E820AAAA80000000000000000000",
INIT_1F => X"AEAAB55007FD74AAAA843DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFF",
INIT_20 => X"2802AA10FFFFFDE0008556AABA5D2ABFFEFFFAAAAAAAF7D57FFEFF7D555555A2",
INIT_21 => X"085542145552ABDFEFFFAA801EFFFFBFDF550000175555504175450055574AAA",
INIT_22 => X"0082A975EF00003DF55555168A00000428AAAAA84021FF007BD54BAAAD17DEBA",
INIT_23 => X"AAFF802ABFF087FFDF5508003FEBA087FD54BA000415400557BD74BAFFD14000",
INIT_24 => X"400AAFBE8ABAF7FFD54AAAAAEA8ABA55557FEAAA2843FF55A2AEA8B55AAAABDE",
INIT_25 => X"00000000000000000000000000000000000000000051554BA002A95555A28417",
INIT_26 => X"C20825D7FE8A92FFFFC70BAE3D155555415178FD7082EAAB550820870BAAA800",
INIT_27 => X"578FFFEBD55557DBEA4AFB550871D7482AA8E3DFFFAAFFD04AA415B52492B6F5",
INIT_28 => X"0E175550051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEFF7A0ADABAEBD",
INIT_29 => X"47BD2482BED57AE921451421555524BDFD7FFA4801D7F7F5FDF55000E1754541",
INIT_2A => X"1C7BD2482E3D1450381C20905EF08003AF55415F6DA38080E2DA82BE8E001EF1",
INIT_2B => X"5BEAAAFB55ABA0BDE02EB8A28BC70075FDF45080A3AEAA007BD24821C0412428",
INIT_2C => X"AA14209557DA28E15400BEF1EFA92FFFFD24BAB6A4A8A82495F78E92AA843DF4",
INIT_2D => X"B450800174BAA680000000000000000000000000000000000000000000055524",
INIT_2E => X"00BA007BC0000FFD542000557FE8A00F3FFD54BAAAD15754508556AB45002AA8",
INIT_2F => X"AABEFFB803DEAAAAD56ABEFAAD5575EFF7803DF45085557410AEAABDFEFAAFBC",
INIT_30 => X"57FF55082E97555002E955550C55554BAFFAEBDE10F7FBFDEBA007BFDE005D2A",
INIT_31 => X"2ABFE00F7AA821FF557FC0010F7D168A105D554214551003FF45FF8400145FFD",
INIT_32 => X"87FC20105504000AA597FC2010A2D1554AA5500021EF000028B55087BFDEBA04",
INIT_33 => X"007FE8A00A2803FF45F7AABDF55AA843FE10AEAAAAB4500557FF55082EA8AAA0",
INIT_34 => X"00000000000055400BA5504155EFAAAE95410F7D57DE00FFFBC00AAFB8028A00",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"A140084000080048040100000202026040000000180800080200010048510204",
INIT_02 => X"080108000090000004655C000080000051000000000402400800000009000010",
INIT_03 => X"0000000100300C40842240000210810002800584488000103080894288800000",
INIT_04 => X"0002584280A2C21000110300100000100220C8C910A032541000090A00643000",
INIT_05 => X"04092A001400D100410A002140004020140001A9005000004810A1C0044D2800",
INIT_06 => X"0360000010EFFD229911C9911820002080258A09A2D3E102137FE0094910A222",
INIT_07 => X"0000004000220400120000090C0810210A040034A040000046180810000C4907",
INIT_08 => X"80404050D88C24510001400042008088090004012000000000010F8102041320",
INIT_09 => X"20080120024030A4090200828C880208002044C0843B44100228A1585C81740A",
INIT_0A => X"142180860A84802042C82180D0010039039390200008B20E2300086800400640",
INIT_0B => X"003000091084190644810502D0A16850B4285B14A688011A1409212008F05E20",
INIT_0C => X"400104080010001E0FF00010000010001E0FF0001002200A1300000000000080",
INIT_0D => X"000080000010001E0FF00010000010001E0FF000100440000040F517CF600000",
INIT_0E => X"E587F9E000004008100800008000ED0FC7E000004000804000000809963F1F80",
INIT_0F => X"36000100202C0020100000000802419660CFE7C0F00000000800810040000040",
INIT_10 => X"0618E7B0000800000003F80FFF0000200018021000030C73D80004000000585F",
INIT_11 => X"078A8FCF600000201802008001006AA3F1F80000400000000B0BD6C000200000",
INIT_12 => X"0041120370DCAD1FC18000000040180200800005D5C3FD800000806008100000",
INIT_13 => X"48A480072284983230101402200200111103202420000880C218000150100800",
INIT_14 => X"2B888A4500048240C08400843204502000890001000415E12480003002944281",
INIT_15 => X"0480004800048000480004800004002240020854884000901212140011C01079",
INIT_16 => X"346D19D1A4C08028904C4E1D7224086590800420044040020004004480004800",
INIT_17 => X"68DA368DA368DA368DA368DA368DA1685A1685A1685A1685A1685A168DA36CDA",
INIT_18 => X"8DA3685A1685A1685A1685A368DA368DA368DA3685A1685A1685A1685A1685A1",
INIT_19 => X"40000000000000000068DA368DA368DA1685A1685A1685A1685A368DA368DA36",
INIT_1A => X"3CF3CF6FE23CCD8D00A281F5B2DB2CA78A543EBC57A10A245DA975D640088884",
INIT_1B => X"3E1F0F87C3E1F0F87CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"5DA9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0F87C",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00B",
INIT_1E => X"40000000043DF55087BC01EF007FD75FFFF84000AAFF80000000000000000000",
INIT_1F => X"2EBFE10A28028AAAAAFBC00AAF7D5575455D557DFEF002AAAB55002E820AAAA8",
INIT_20 => X"2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFAA95545552ABFE00087BC00AA08",
INIT_21 => X"007FD74AAAAD57FF45002A975FF007BE8BFFA2FBFFFFFAAD5400AAFF843DFEFA",
INIT_22 => X"5AAFBE8A00082A97410F7D5555EFAAAAAAAAAF7D57FFEFF7D555555A2AEAAB55",
INIT_23 => X"450055574AAA2802AA10FFFFFDE0008556AABA5D2ABFFEFFFAA8200055555554",
INIT_24 => X"F55000017555550417545000015545087BC2010AAD54014500516ABFFA2AABDF",
INIT_25 => X"0000000000000000000000000000000000000000002ABDFEFFFAA801EFFFFBFD",
INIT_26 => X"AAB550820870BAAA8407000140038F450075C71FF087BD75D7FF84050BAEB800",
INIT_27 => X"AB8E10007FC50BA002ABFE00AA8A2AABABEFFC70BAE3D155555415178FD7082E",
INIT_28 => X"DB45082EB8E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92FFA497545552",
INIT_29 => X"BD55557DBEA4AFB550871D7482AAD17DF451C24955EF0875EFBD7B6F1FFFC7BE",
INIT_2A => X"F7AA87000415B5057DAAFBE8A10082092410EBD5505EFB6A0ADABAEBD578FFFE",
INIT_2B => X"D005B6ABC7B6AABFFED0051574BAB68A2DA00FFFFFFE38085F6FA92552AB8FEF",
INIT_2C => X"D7FFA4801D7F7F5FDF55000E17545410E17555000E17545007BC0000BED14217",
INIT_2D => X"555F784174AAA280000000000000000000000000000000000000000000024BDF",
INIT_2E => X"754508556AB45002AA8B450800174BAA684174105D042AB550055555FF007BD7",
INIT_2F => X"E8A00F384175555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7FFD54BAAAD15",
INIT_30 => X"57DF55FFD57DF55FFFBD5400A2AABDFEFAAFBC00BA007BC0000FFD542000557F",
INIT_31 => X"803DEAAAAD56ABEFAAD5575EFF7803DF45085557410AED17FF455D04155FF005",
INIT_32 => X"07BFDE005D2AAABEFFBAE97410087BC21EFA2FFEAA00000002010A2D5421FFFF",
INIT_33 => X"087BC0010FFD1401EF087FE8B55FFAEBDFEF0855554BAFFAEBDE10F7FBFDEBA0",
INIT_34 => X"000000000000003FF45FF8400145FFD57FF55082E97555002E955550C2E95555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000002000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000006",
INIT_01 => X"0000098218302849180060000C004260413C0A61590001D90213C80000110200",
INIT_02 => X"680108220010000054400C00008000004100000001200240080080000908A011",
INIT_03 => X"000A0000040020400002021000000008428065044880001030818C0008C10000",
INIT_04 => X"00005042882A8210003000000800001000806080100040140080040800003140",
INIT_05 => X"0400000840000098410800010001002000000000004000002010000040002000",
INIT_06 => X"03600810100001220911E0911902000020200200A253E8000C0010080800004C",
INIT_07 => X"000408C0002204400200000B080000010C040004A0400000C0000810000C5901",
INIT_08 => X"000008002A84300000014000C2008088090008002000000000030F8000001220",
INIT_09 => X"0008012100000200001200820888010800200000000840100028800004801440",
INIT_0A => X"000090220000040400480000D0010009049090200008B2022384800802010000",
INIT_0B => X"001000090001090A4C81240050A328519428CA14328C840A5820000101500400",
INIT_0C => X"00510008100400000000A00000100400000000A00000000A12000000000000B0",
INIT_0D => X"00012000100080000000A00000100080000000A0000540000000000000000000",
INIT_0E => X"00000000000000A8000900010000000000000000060000420004000000000000",
INIT_0F => X"0000024000240000102000000080000000000000000000240000800140000000",
INIT_10 => X"0080000000120CFC000000000000000001280013E010000000000900F8040000",
INIT_11 => X"2000000000000001480006D5801000000000000000091F0000800000004807C0",
INIT_12 => X"901A800080000000000000000820080006DD000000000000000002A00019DC00",
INIT_13 => X"0200800522C01252501086222082000010012024200000048019502000000C32",
INIT_14 => X"0080004501000200089400005200D0820008000000104C4800010600BC228404",
INIT_15 => X"0001040010000104001000010440080000822900000000801010500A13404111",
INIT_16 => X"32851951A0CA8080924C06403600086491900224002200400440104001040010",
INIT_17 => X"284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A128CA328CA",
INIT_18 => X"84A1284A1284A1284A1284A328CA328CA328CA328CA328CA328CA328CA328CA3",
INIT_19 => X"10000000000000000028CA328CA328CA328CA328CA328CA328CA1284A1284A12",
INIT_1A => X"69A69A250B61004055CD1439248209070CCCF48DE68A8900401038E2550A0010",
INIT_1B => X"341A0D068341A0D068A28A28A28A28A28A28A28A28A28A28A28A28A29A69A69A",
INIT_1C => X"56C1A0D269341A0D068349A4D068349A4D068341A0D269341A0D269341A0D068",
INIT_1D => X"0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE052",
INIT_1E => X"57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D00000000000000000000",
INIT_1F => X"D1575EF00557DF555D040000000043DF55087BC01EF007FD75FFFF84000AAFFD",
INIT_20 => X"7D5575455D557DFEF002AAAB55002E820AAAA843DFEF00517DEBA007BFDFEFFF",
INIT_21 => X"A28028AAAAAAABDF45F7803FFEF555568AAAF7802AA00FFFBD7555087BC00AAF",
INIT_22 => X"5087BD54BA550417400085155555082A95545552ABFE00087BC00AA082EBFE10",
INIT_23 => X"555D043DFEFA2FBD54BA5555554BAAAFBC20BA5D7BEAAAAFFFBC00AA552E9554",
INIT_24 => X"BFFA2FBFFFFFAAD5400AAFF8402000A2FFFDF555D7BE8BFF5D51575EFA280175",
INIT_25 => X"000000000000000000000000000000000000000000557FF45002A975FF007BE8",
INIT_26 => X"D75D7FF84050BAEBDF78F45B68010482415B471C7E3DF451EFBEFBFAF4549000",
INIT_27 => X"17DE82007FFAFEFE3DB505EF1C5B7AF45490407000140038F450075C71FF087B",
INIT_28 => X"FFD55451C7FC70BAE3D155555415178FD7082EAAB550820870BAAA8438FFF005",
INIT_29 => X"07FC50BA002ABFE00AA8A2AABABEAEB8F45F78A3DFD741516DAAAE38E2DA28EB",
INIT_2A => X"FFFFC20BA5D2E905550071D54825D0A1543808515756D1C2497545552AB8E100",
INIT_2B => X"F5D55505FFBE801256D490E3DFFFAAFFD04AA415B52492B6F5C20825D7FE8A92",
INIT_2C => X"451C24955EF0875EFBD7B6F1FFFC7BEDB45082EB8002000AAFFFDF6D417FEABE",
INIT_2D => X"5EFF7FBE8B5500000000000000000000000000000000000000000000000517DF",
INIT_2E => X"AB550055555FF007BD7555F784174AAA2FBEAB45F78402010007BD5545AAFFD5",
INIT_2F => X"174BAA68028BEF00517FE10007BE8BFFAAFFC01FF557FE8B550004174105D042",
INIT_30 => X"57FEAAAAAEBFEAAAAFFD5545557FD54BAAAD15754508556AB45002AA8B450800",
INIT_31 => X"04175555D2EA8A00087BD74BA082EBDE10AAAEA8ABAF7AAAAB45F7AEBFF45085",
INIT_32 => X"FD542000557FE8A00F3FFC00BA552E80145005557400552A954BA0051575EF55",
INIT_33 => X"A2FBFDFFF007FE8BFF5551401EFF784021FF002ABDFEFAAFBC00BA007BC0000F",
INIT_34 => X"000000000000517FF455D04155FF00557DF55FFD57DF55FFFBD5400A28400010",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000004000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A14009801830084C182060000C10424840000000080000080200000000110204",
INIT_02 => X"0801080200100000046558040080000041000000002402400800000009008010",
INIT_03 => X"00020201040000D0842242024210810802006400088000003080054288C10000",
INIT_04 => X"0000400088020000003020002000001002A0E881108032100002000800203040",
INIT_05 => X"04092A081000411841480001000000201000012800400010001081C040402000",
INIT_06 => X"03600810100001220001E0001802002020240208000369001500100909000266",
INIT_07 => X"0000004000220440020000090C0810210A040004A0410000C0000810000C4901",
INIT_08 => X"0040480000802100100140004200808809000C002000000000010F8102041320",
INIT_09 => X"2008012000000000000200828888800808000410800840100220211850004442",
INIT_0A => X"040180240A80800442400004C0010000060210200008B2022304880800010000",
INIT_0B => X"0030000000010008008020020100008000400120800004004821202001A05A00",
INIT_0C => X"40510008101480000000A01004101480000000A0100000001300410402080080",
INIT_0D => X"0001A004101480000000A01004101480000000A0100540000040000000000000",
INIT_0E => X"00000000000040A8000900018040000000000000460800420004090000000000",
INIT_0F => X"0000034000082000102000000080028000000000000000240800800140000040",
INIT_10 => X"20900000001A00000002000000000020013000100010480000000D0000040440",
INIT_11 => X"2018000000000021500000800010440000000000400900008088000000680000",
INIT_12 => X"000000008200800000000000086010000080000100000000000082C000100000",
INIT_13 => X"000080000004924040008020000200101100004000000000C019500050000800",
INIT_14 => X"2B088A4541008240001000804000108280800001001051A12481041080801010",
INIT_15 => X"4480004800048004480044800044000240022100884000901210440003C14110",
INIT_16 => X"06E00000044200009849485D4020080000140004046240020044000480044800",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802000000400",
INIT_18 => X"0000000000000000000000020080200802008020080200802008020080200802",
INIT_19 => X"1000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"1451451AA654199951A24454514514F0CA940FE0D39712615FAD555204428290",
INIT_1B => X"CA6532994CA65329945145145145145145145145145145145145145145145145",
INIT_1C => X"670E572994CA6532994CAE572B95CA6532994CA6532B95CAE572994CA6532994",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE01C",
INIT_1E => X"03FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF0800000000000000000000",
INIT_1F => X"7FFDF45FFFBC2010AAD57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D0",
INIT_20 => X"0043DF55087BC01EF007FD75FFFF84000AAFF8002155AAFFE8B45AAD54000008",
INIT_21 => X"00557DF555D517FEBA082A801EFF7FBD5400FFD568B555D00155EF0804000000",
INIT_22 => X"AF7FBFDE00A2FBC0145005168A10AA843DFEF00517DEBA007BFDFEFFFD1575EF",
INIT_23 => X"EF5D7BC00AAF7D5575455D557DFEF002AAAB55002E820AAAA803FEBA082AAAAA",
INIT_24 => X"AAAF7802AA00FFFBD7555082E82155FFAEAAB55AAD568B455D00154BAFFFBD75",
INIT_25 => X"0000000000000000000000000000000000000000002ABDF45F7803FFEF555568",
INIT_26 => X"451EFBEFBFAF4549003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC700000",
INIT_27 => X"5EDB6DAADF470280075FFF45E3F1C7038A2DF78F45B68010482415B471C7E3DF",
INIT_28 => X"0A175C7000407000140038F450075C71FF087BD75D7FF84050BAEB8002155BEF",
INIT_29 => X"07FFAFEFE3DB505EF1C5B7AF45495B7DEAA0824851EFEBFBD2410EBD168B7D41",
INIT_2A => X"AA8038EAA0824A8AAAEBF5FAE28AAF1C2155005F68A10A28438FFF00517DE820",
INIT_2B => X"D4104104AAF7F1D75EF557FC70BAE3D155555415178FD7082EAAB550820870BA",
INIT_2C => X"45F78A3DFD741516DAAAE38E2DA28EBFFD55451C2087155EBA4A8B7DAADF68B7",
INIT_2D => X"FEFA2AEAAB55000000000000000000000000000000000000000000000002EB8F",
INIT_2E => X"2010007BD5545AAFFD55EFF7FBE8B5500043FE00F7D17FEBAA2D5574BAAAD17D",
INIT_2F => X"174AAA28002155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAB45F7840",
INIT_30 => X"BC2000AAD16ABFF002A975450004174105D042AB550055555FF007BD7555F784",
INIT_31 => X"8028BEF00517FE10007BE8BFFAAFFC01FF557FE8B55007FFDEAA0004175FFA2F",
INIT_32 => X"02AA8B450800174BAA68428AAA08042AABAAAD56AABAAAD140155087FEAA10A2",
INIT_33 => X"A2842ABEFAAFBE8BFF0004020AAFFD5555EF557FD54BAAAD15754508556AB450",
INIT_34 => X"0000000000002AAAB45F7AEBFF4508557FEAAAAAEBFEAAAAFFD5545550015555",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000047FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B83008481800E0000C26426040000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"00080D4912E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"000048048002400048150000000002504230C899109032100020160880223000",
INIT_05 => X"040B2A229100410041088011100022201200012840440000B01088C0005C2400",
INIT_06 => X"03286A287E4003225021C5021880C02000A40249048363A5990010090908022A",
INIT_07 => X"8320694044222987020C80152D8910210A0400252B74200045C86810000C5B05",
INIT_08 => X"00404126509804400501400242C0B0B83B0134702000000000191FA162841324",
INIT_09 => X"2008013002000220001240820F8B2A08000040409018401001200159D80D64AA",
INIT_0A => X"91019B02080885200042E098C00101B0070310200008B60A23A51B2802067327",
INIT_0B => X"003000080802500C088325828102408120409120940680100504022148504440",
INIT_0C => X"1501D5761B011986695014A96E1A8119865A5018C5A0A00012004104020808B0",
INIT_0D => X"A2600AAE1A811986695014A96E1B0119865A5018C5AF0062C38A4DB680A0D824",
INIT_0E => X"1DB528802CAB184E8F4101621B1BAC845542056A289A1BB2078A922DA2A8B180",
INIT_0F => X"7A3D94392000224ACDE215883078681B5C05AA429189B60AC43CEC7F0272C384",
INIT_10 => X"134CD551BCA1C90006C0C2958502861120C003104289A668B8CAB27010633831",
INIT_11 => X"82806CA64090B89E015AAA880E48382EB8804B020A06020C67061BC785938085",
INIT_12 => X"470126C6284B2D20410AB4503089C00A8280819A5539D503336D61056ABA0062",
INIT_13 => X"000080060040142020015001004A00080042004000E8089C9003066E03513E41",
INIT_14 => X"010CBA45367082014000908020349320008000A1000C09A9348498B000000000",
INIT_15 => X"C32A0832A0C32A0C32A0832A0C19504195040040000000801010028001400010",
INIT_16 => X"2468118104400000904C0C0964200841010954000444D280140050C32A0832A0",
INIT_17 => X"4090240902409024090240902409024090240902409024090240902409024090",
INIT_18 => X"0100401004010040100401024090240902409024090240902409024090240902",
INIT_19 => X"0000000000000000004010040100401004010040100401004010040100401004",
INIT_1A => X"410410502A441495418984700000005088804180C0B10A04D0A7104201400284",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000010410410",
INIT_1C => X"7800000000000000201000000000000000000008040000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE060",
INIT_1E => X"4155EFAA842ABEFA280155EFFFFBC01EF0855400005500000000000000000000",
INIT_1F => X"FBFFF4508514000000003FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF080",
INIT_20 => X"280154BA5555401EFFFD5421EFA2FFFFF555D51575FFA2FFD75FF550015400FF",
INIT_21 => X"FFFBC2010AAD568AAAAAD142145FF80155EF0051555FF0804155FFF7D57DF45A",
INIT_22 => X"008001540008514215555003DFFFA28002155AAFFE8B45AAD540000087FFDF45",
INIT_23 => X"0000040000000043DF55087BC01EF007FD75FFFF84000AAFF802ABFFA2AABFE1",
INIT_24 => X"400FFD568B555D00155EF085168B45085142010FFAE800AA5D7BFDF45F7FFEAA",
INIT_25 => X"000000000000000000000000000000000000000000517FEBA082A801EFF7FBD5",
INIT_26 => X"7DF7DA2AEB8FC70000175EFB6802DBC7BE8A155EFE3FBC71FF145B4203855000",
INIT_27 => X"5D05EF550E15400E3F1FFF7D085B420381C003DE10BEF5EDAAAAAD547038EBD5",
INIT_28 => X"04105C7F7DF78F45B68010482415B471C7E3DF451EFBEFBFAF45495F575FFBEF",
INIT_29 => X"ADF470280075FFF45E3F1C7038A2DB68ABAB6D145145FF84155D7085B555C714",
INIT_2A => X"EB8428BEFBEA4BDE28140A1543800514515549003FFC7BE8002155BEF5EDB6DA",
INIT_2B => X"2417FFFF7DE3F1EFA10140407000140038F450075C71FF087BD75D7FF84050BA",
INIT_2C => X"AA0824851EFEBFBD2410EBD168B7D410A175C7005B6DB55145140000FFAE8508",
INIT_2D => X"5EF557BC20AA5D0000000000000000000000000000000000000000000005B7DE",
INIT_2E => X"FEBAA2D5574BAAAD17DFEFA2AEAAB550004175FFF7803DF45FFAE955EFAAFBD5",
INIT_2F => X"E8B55007FD75FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D043FE00F7D17",
INIT_30 => X"015555007FD5545550400145FFFBEAB45F78402010007BD5545AAFFD55EFF7FB",
INIT_31 => X"8002155FFD17FFFFA2FBD74BA00557FF45A2D5554AAA2FBEAAAAFFD555545FF8",
INIT_32 => X"07BD7555F784174AAA2842ABEFFF803DEAA5D2E974AA00515754500003FF55FF",
INIT_33 => X"555540000FFAE97410007BFFFFFA2D57FE105D04174105D042AB550055555FF0",
INIT_34 => X"0000000000007FFDEAA0004175FFA2FBC2000AAD16ABFF002A97545007FFFF45",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000004000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C048000C048400380000007024040000000080000088200002802153231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"421A0A0012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"02004000890200001837800001998C31C090609C104000102002140900003548",
INIT_05 => X"0402002BC200009841090001200006200800000020480010A4100100001C2000",
INIT_06 => X"033432287FC003230001D0001806C0060CB0622000037085C800100C0C200008",
INIT_07 => X"135038CE64B663DFA314C803292140890C0601F472D1640051F80C10020C493F",
INIT_08 => X"00000167C081000011814004C20481A92940EA7A3020480000071F846890162E",
INIT_09 => X"D40C01240008000080024082488BAF08000020000208401004300421800F04F8",
INIT_0A => X"F9F80FA0200E0BF40063FF9DC0010000180018200408B27E234913E900067F04",
INIT_0B => X"001100002002801000A04200000000000000000000029D204B7C0382FD0100F3",
INIT_0C => X"9628F97E0B348EDAC3900F6EFA0B158EDA93900F6EE230381208008001007A80",
INIT_0D => X"EAE64BCA0B158EDAC3900F6EFA0B348EDA93900F6EE8421392C96B1237E0D8BD",
INIT_0E => X"4CAEAD412EDD2B47CFF812A383430C669E622DBC31D73F6006A5891533EF9500",
INIT_0F => X"2E19B8BA30E022DAD8C100CA39E8CEBE66C2B083798D341B10DE7E14400392C7",
INIT_10 => X"32966471A9C5DD00B12728D5360234D62A49FAB442994B3238D4E2FB10463665",
INIT_11 => X"F0FABAC800DA550C29F36A8A2554E48A6430469392526208C6CC95C33717D885",
INIT_12 => X"2B416A51B60585A5C28895962502E9F36A828C4999AF580395542D27CDBA0020",
INIT_13 => X"0000800000001E404011F066000A000EE040000000873FB80B8A00EF03F56CC1",
INIT_14 => X"2284304D667C06CC6816B300403C13E2000000460010400000010CE080801010",
INIT_15 => X"872F0872F0C72F0872F0872F0C597863978421000800209010104ACA03414110",
INIT_16 => X"01000000104280009048004000000800001D5E05182493C5BC5AF0872F0C72F0",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0802008020080200802008000000000000000000000000000000000000000000",
INIT_19 => X"1000000000000000000080200802008020080200802008020080200802008020",
INIT_1A => X"492492240F010000146E502D4514510246088881360A95118B120CB054420210",
INIT_1B => X"6432190C86432190C82082082082082082082082082082082082082092492492",
INIT_1C => X"7FEB2592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2590C8",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"5421FF00042ABEFFF8400010082EAABFF55002ABEF0800000000000000000000",
INIT_1F => X"002ABEFFFFBD54000004155EFAA842ABEFA280155EFFFFBC01EF085540000555",
INIT_20 => X"AFBE8AAAA2D540000F7D57DF55A2AABFFEF08556AA10000028AAAFFD15541000",
INIT_21 => X"085140000005168AAA087BFFFFF5D04001FF00041554555557FE005D003FE10A",
INIT_22 => X"F0851555FF082AA8B55F7AEA8BEF5551575FFA2FFD75FF550015400FFFBFFF45",
INIT_23 => X"10AAD57DF45A280154BA5555401EFFFD5421EFA2FFFFF555D0000145082E955F",
INIT_24 => X"5EF0051555FF0804155FFF7842AA100000020BAAA801541055042ABEFFFFBD54",
INIT_25 => X"0000000000000000000000000000000000000000005568AAAAAD142145FF8015",
INIT_26 => X"C71FF145B42038555F401D71C0A2DBC7EB80000280824ADBD7490E28BEF08000",
INIT_27 => X"A2DA82FFDB5243800002FBD7EBFBD24101C00175EFB6802DBC7BE8A155EFE3FB",
INIT_28 => X"5B7AE1041003DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7005F6AA381C0",
INIT_29 => X"50E15400E3F1FFF7D085B420381C5B6AA82147FF8FEF410E001FF000E1755555",
INIT_2A => X"49000017D142E905EF1451525C7082AADB45F7AEA8BEF555F575FFBEF5D05EF5",
INIT_2B => X"041002FBEFEBFBD2410AADF78F45B68010482415B471C7E3DF451EFBEFBFAF45",
INIT_2C => X"BAB6D145145FF84155D7085B555C71404105C7F7842FA381C0A00082AA8A1041",
INIT_2D => X"F55002AA8BEF000000000000000000000000000000000000000000000005B68A",
INIT_2E => X"DF45FFAE955EFAAFBD55EF557BC20AA5D7BC01555D2EBFF55A284000AA08003F",
INIT_2F => X"AAB55007BE8AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D04175FFF7803",
INIT_30 => X"E821FF082A97555557FE8A0000043FE00F7D17FEBAA2D5574BAAAD17DFEFA2AE",
INIT_31 => X"7FD75FFF7D5401EF5D2E97410AAD17DFEF007FC20AA5D7BE8A005D7FEABFF002",
INIT_32 => X"AFFD55EFF7FBE8B550004001FF5D2A801EF5D5142145082EBFF55F7AAAABEF5D",
INIT_33 => X"552A82010A2AA8000008043FFFFA2FBC2010A2FBEAB45F78402010007BD5545A",
INIT_34 => X"0000000000007BEAAAAFFD555545FF8015555007FD5545550400145FF843DEAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400986B830E84D182260000C1042684001000008220008A20019080A510200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00020201926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"00104884880A4400403003005800027102A0E8C110D83210642EA809C0203040",
INIT_05 => X"04092A08138041184109C001380000201A008128044E00754010C9C192D82400",
INIT_06 => X"032C7E201800012372A1D72A180000204024024954A3670819001009092C0222",
INIT_07 => X"0164004000220B40020C80052C0A12292A040005715540015E006810001C4B01",
INIT_08 => X"0040549032881001140140024200808839005C002010800000155F8122851320",
INIT_09 => X"6008012C80481284881280825A988008000040808629441005B3071859006442",
INIT_0A => X"0001B0200810940400720005C0030192072310200028B6022346080802E001A5",
INIT_0B => X"003000206822F20CA8826AC2A14250A128509528954404144C20042501004000",
INIT_0C => X"03D404A41AA5B7344C10B383081BA4B7341C10B3831034081200000000000430",
INIT_0D => X"5A2B2C381BA4B7344C10B383081AA5B7341C10B383110218CB0E54C2EA404A4F",
INIT_0E => X"3548B3A008E730A01AB113A5524E6ACA678001CE3E20A5B284ED1132909C7288",
INIT_0F => X"0A3C066430202021252991C22C99731014AC3CC0C0B8182597A801610218CB0C",
INIT_10 => X"A5C8825194332B018A444AEA2701288A15A151EC5952E44128CA194517354C18",
INIT_11 => X"635232D50048A411C158BB0A7910142C771804C8A0ADA2E6A983014780CA28B2",
INIT_12 => X"6E4023F8BE8E3E1E0109472C3EB50158BB02D09852745F80112C428562EE0353",
INIT_13 => X"00008002414032646000826080C20001104240480068001C9B9150A000029704",
INIT_14 => X"1118BA4510008241C80290882400908000A000A1000809A93485D61000000000",
INIT_15 => X"40000000000000040000000000000020000000040000008010122A8201410058",
INIT_16 => X"246A10A1044101A89A4D0C096420184321040002844840000000004000000000",
INIT_17 => X"5094250942509425094250942509425094250942509425094250942509425094",
INIT_18 => X"0942509425094250942509425094250942509425094250942509425094250942",
INIT_19 => X"0000000000000000005094250942509425094250942509425094250942509425",
INIT_1A => X"75D75D7FEDFDFDFDFBEEF9DD555555F7EEFF3F7DF7FF3E7E1FBF7DF7E24502A8",
INIT_1B => X"FAFD7EBF5FAFD7EBF5D75D75D75D75D75D75D75D75D75D75D75D75D75D75D75D",
INIT_1C => X"7FEFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F780000000000000000000",
INIT_1F => X"AA97400AAD540155A2D5421FF00042ABEFFF8400010082EAABFF55002ABEF085",
INIT_20 => X"A842ABEFA280155EFFFFBC01EF08554000055043DEBAF7843FFFFF7AABDF55A2",
INIT_21 => X"FFFBD5400005568A1055043DEBAAAFFE8B45557FD7410552EAAABAAA84155EFA",
INIT_22 => X"AA2FFE8ABAAA8428A00087BD7555FFD56AA10000028AAAFFD15541000002ABEF",
INIT_23 => X"55A2803FE10AAFBE8AAAA2D540000F7D57DF55A2AABFFEF085557545FFD17DEB",
INIT_24 => X"1FF00041554555557FE005D0000155557BEAABA5D2ABDF450851420AA5D7FD55",
INIT_25 => X"0000000000000000000000000000000000000000005168AAA087BFFFFF5D0400",
INIT_26 => X"ADBD7490E28BEF08516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EB800",
INIT_27 => X"03FFD7EBA4BDF45AAAA90410BEDF45155A2DF401D71C0A2DBC7EB80000280824",
INIT_28 => X"2AAFA82B680175EFB6802DBC7BE8A155EFE3FBC71FF145B42038550E38E92EB8",
INIT_29 => X"FDB5243800002FBD7EBFBD24101C556FA38490A3FE92BEFFEAB45417FD24385D",
INIT_2A => X"00515056DE3D17FE92BEF1EFA92AA8428A10007FD557DFFDF6AA381C0A2DA82F",
INIT_2B => X"5085B400925D7FD557DA2803DE10BEF5EDAAAAAD547038EBD57DF7DA2AEB8FC7",
INIT_2C => X"82147FF8FEF410E001FF000E17555555B7AE10410E00155497FEFABA4120B8F5",
INIT_2D => X"ABAA2FBD7545AA8000000000000000000000000000000000000000000005B6AA",
INIT_2E => X"FF55A284000AA08003FF55002AA8BEF00517FE00082EBDF45AA8428A10085568",
INIT_2F => X"C20AA5D2EA8A00A2803DF45AA843DF55AAAE82000F7FBD5545AAFBC01555D2EB",
INIT_30 => X"FE8B55087FC00BA552ABFE10F784175FFF7803DF45FFAE955EFAAFBD55EF557B",
INIT_31 => X"FBE8AAA5D2EBDE00FFFFC00AA08003FF55A2FBC00105D517FEAA082EBFE10F7F",
INIT_32 => X"AD17DFEFA2AEAAB550051401FFA2D57FE10F7D57DE00AA842AA00007FD75FFF7",
INIT_33 => X"007BFDEAA08042AB45087FC0010557FD55FFAA843FE00F7D17FEBAA2D5574BAA",
INIT_34 => X"0000000000007BE8A005D7FEABFF002E821FF082A97555557FE8A00002E82155",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000067FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"0002074F200904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000480488024000403000000000001002A0E881108032100002000800203040",
INIT_05 => X"04092A081000411841080001000000201000012800400010001081C000402000",
INIT_06 => X"033D7880500001221021C1021800002000240249048361001100100909000222",
INIT_07 => X"9020304000220050020480152D0A142D0A8400043B45400040006810000C5901",
INIT_08 => X"0040400010880000100140024280808829029C002000000000053FA142051324",
INIT_09 => X"6008012000000000000200820888800800004000800840100020011858006442",
INIT_0A => X"000110200800840400400005C0010190070310200008B202236D080802000001",
INIT_0B => X"003000000000100C088020028102408120409120940404104C20002101004000",
INIT_0C => X"2050805210040000B0E0A0000210040000E0E0A0000190081200000000000000",
INIT_0D => X"0111300210008000B0E0A0000210008000E0E0A0000B02740421A0E5D1A02400",
INIT_0E => X"C0715C40110080A4006110510C14D18178E01200860008920106460D4501CB00",
INIT_0F => X"500002411420220080220C0093C38923240ABBC00905C33C6000400F02740412",
INIT_10 => X"9682398000120800658992F3C700C3018120000041DB011CC000090012565306",
INIT_11 => X"B7A0B1E240240A8340000200067EAA8CB65809240C09024A4AE0CA0000480083",
INIT_12 => X"00845C7DB0D0200900422ACA4B28000002002B46867DBC002A830280000800F7",
INIT_13 => X"000080020040126060008020000200000042004005800004801150A003412440",
INIT_14 => X"01088A4500008240000000802000908000800001000009A92481041000000000",
INIT_15 => X"0000000000400000000000000400000000000000000000801010000001410010",
INIT_16 => X"246810810440000090480C096420084101040000044040000000004000040000",
INIT_17 => X"4090240902409024090240902409024090240902409024090240902409024090",
INIT_18 => X"0902409024090240902409024090240902409024090240902409024090240902",
INIT_19 => X"0000000000000000004090240902409024090240902409024090240902409024",
INIT_1A => X"3CF3CF3FE77DDDDD55E6D5FCF3CF3DF7CE5C8FF0F7BE9D75CF9F7DF650400280",
INIT_1B => X"FE7F3F9FCFE7F3F9FCF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"8007F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE07F",
INIT_1E => X"17DF45AAD157400007BEAAAAAAAE955555D5568A105D00000000000000000000",
INIT_1F => X"AA800AAF784020AAF7D56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7D",
INIT_20 => X"0042ABEFFF8400010082EAABFF55002ABEF085155400FFD1420100055574AAA2",
INIT_21 => X"AAD540155A28028B550051574005D7FFFE105D7BD7545A284020BA0055421FF0",
INIT_22 => X"00851421FF5D7FFDEBA085168B45FF843DEBAF7843FFFFF7AABDF55A2AA97400",
INIT_23 => X"FF5504155EFAA842ABEFA280155EFFFFBC01EF08554000055002AB455D514201",
INIT_24 => X"B45557FD7410552EAAABAAA8017400AAD140000002EBFFEFA2AAA8BEFF780021",
INIT_25 => X"0000000000000000000000000000000000000000005568A1055043DEBAAAFFE8",
INIT_26 => X"F8E38E3DF45155EBD17FF6DAADB504001C71EDA82AAA0955455D556DA0049000",
INIT_27 => X"B420101C55554AAAAA480082FF84000BAEBD16DA82410A3FFD7AAA4B8E824971",
INIT_28 => X"8405092085F401D71C0A2DBC7EB80000280824ADBD7490E28BEF085157428FFD",
INIT_29 => X"BA4BDF45AAAA90410BEDF45155A28E2AB7D0051504005D71F8E004975D556DB6",
INIT_2A => X"550028B6D5D51420101C5B401EF417BFAEAA08516AB45E38E38E92EB803FFD7E",
INIT_2B => X"7A2AEAFBC7EB80071FF5500175EFB6802DBC7BE8A155EFE3FBC71FF145B42038",
INIT_2C => X"38490A3FE92BEFFEAB45417FD24385D2AAFA82B68015400AADB40000082EBFFC",
INIT_2D => X"54555557FE1000000000000000000000000000000000000000000000000556FA",
INIT_2E => X"DF45AA8428A10085568ABAA2FBD7545AAD17DFFFAAFFC200055557DE00A28015",
INIT_2F => X"A8BEF0051554AAFFFFC00105D55554BAA28400000F784020BAAAD17FE00082EB",
INIT_30 => X"568A000051575FFF78415410087BC01555D2EBFF55A284000AA08003FF55002A",
INIT_31 => X"AEA8A00A2803DF45AA843DF55AAAE82000F7FBD5545AAAEAABFF0051400105D5",
INIT_32 => X"AFBD55EF557BC20AA5D042ABFF555142000557FC01EF007FEAABA00556AB55A2",
INIT_33 => X"A2FBC0010082EBDF55A2AABDF45A284175FF5D04175FFF7803DF45FFAE955EFA",
INIT_34 => X"000000000000517FEAA082EBFE10F7FFE8B55087FC00BA552ABFE10F78415400",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000100000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"000440009282000001100000000000100220C8811080321000000228002A3000",
INIT_05 => X"04092A0010004300418800510000A6201000012A64400000145080C000422000",
INIT_06 => X"032B1800100001220001C00018821020402402080003772019001009090002AA",
INIT_07 => X"0000004000220000021840010C8912250A0400042044400040006810000C4901",
INIT_08 => X"0040400022810000058140024280A0A8190004002030C00000016F8122041320",
INIT_09 => X"E0080120000000000002C0820888008800000000800840100020011850004402",
INIT_0A => X"00013000080094000062000180010180060210200008B2022304080800000003",
INIT_0B => X"0030000000000008008020020000000000000100800000000000002500004000",
INIT_0C => X"0000000010108000000000000010108000000000000230001200000000000420",
INIT_0D => X"0000000010140000000000000010140000000000000100000040000000000000",
INIT_0E => X"0000000000000000000100008040000000000000000000020000090000000000",
INIT_0F => X"0000000030002000406000000000068409014000000000000000000100000040",
INIT_10 => X"2010000000000800000201000800000000000000400048000000000010000440",
INIT_11 => X"00184400A0000000000002000000441108800000000002008008000000000080",
INIT_12 => X"0000000242038B82800000000000000002000001000000000000000000080000",
INIT_13 => X"000080000000100000000005C04A000000400000000000000001062000000400",
INIT_14 => X"01088A4500008200000000800000100000800001000001A12480001000000000",
INIT_15 => X"4000040000000000000000000400002000020000000000801010000041400010",
INIT_16 => X"0460000004400000904808094020080000000000044040000000004000040000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000400280",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FC00000804154AA5D00001EFF78428AAA007BC2145F780000000000000000000",
INIT_1F => X"55400AA007FC2000F7D17DF45AAD157400007BEAAAAAAAE955555D5568A105D7",
INIT_20 => X"D043FFFFAAAABDEAA557BFDE00FFD140155F7FBD74AAAAD17DF45F7D1421EF00",
INIT_21 => X"F784020AAF7FFFDF45FF84000BA552ABDFEF08517DF55A2FBEAB555D556AAAA5",
INIT_22 => X"5AAFFEAB45F7843FF45082A801FF005155400FFD1420100055574AAA2AA800AA",
INIT_23 => X"AAA2D5421FF00042ABEFFF8400010082EAABFF55002ABEF087BE8ABA555168B5",
INIT_24 => X"E105D7BD7545A284020BA007FFFE10A284000AA0055401550055574005D2E800",
INIT_25 => X"0000000000000000000000000000000000000000000028B550051574005D7FFF",
INIT_26 => X"955455D556DA004971C7038140012482550E021C7EB8028A821C7BC516DFF800",
INIT_27 => X"17FF45E3DF471C70851400BA0071C5028FFD17FF6DAADB504001C71EDA82AAA0",
INIT_28 => X"FBE8B555D516DA82410A3FFD7AAA4B8E824971F8E38E3DF45155EBF1D5492BED",
INIT_29 => X"C55554AAAAA480082FF84000BAEBF1FFF7DEB8000092552ABFFEF08517DF6DB6",
INIT_2A => X"087FEFA8241516DB55A2FFEAB6DEB843DF551C20801C71C5157428FFDB420101",
INIT_2B => X"5085550428412A85082BEDF401D71C0A2DBC7EB80000280824ADBD7490E28BEF",
INIT_2C => X"7D0051504005D71F8E004975D556DB68405092087FF8E00BE8A02082005F4714",
INIT_2D => X"A00557BD75EFF78000000000000000000000000000000000000000000000E2AB",
INIT_2E => X"200055557DE00A2801554555557FE100055554BA5504000105D2A80145AA842A",
INIT_2F => X"D7545AAD557410F7D57DF55AAFBD55450055420BA0055574BAF7D17DFFFAAFFC",
INIT_30 => X"ABDFFF08517FFFFF7FBEAB455D517FE00082EBDF45AA8428A10085568ABAA2FB",
INIT_31 => X"51554AAFFFFC00105D55554BAA28400000F784020BAAAD57FFEFA28402010552",
INIT_32 => X"8003FF55002AA8BEF007FFDE1000557DF45AAFBE8BEFA2803FF4555040015555",
INIT_33 => X"F7AE80000087BD55450855400BA002A95400F7FBC01555D2EBFF55A284000AA0",
INIT_34 => X"0000000000002EAABFF0051400105D5568A000051575FFF78415410087FEAA10",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000006000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"0202115002BB10080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"2FE962000017102918900948514522CE09200C0D590569398ADBF8CC1E50E480",
INIT_05 => X"5E6023002834854AE41C1E8782F508F2A15B71D412E0AFD9C2990DA56FF0B55A",
INIT_06 => X"82A803B9B9E55402000340003200220A86012D0000000480D02A7960540180A0",
INIT_07 => X"01380C40D890101DBD400901442800817C2901F400868554DE240000A80090CE",
INIT_08 => X"18A9050122004000005665510320C9C90510025A8A00000A0A048F550A440E00",
INIT_09 => X"2A8A562060410280081116C8204D016CB2CB2900080082795804112890000001",
INIT_0A => X"4052E400008176802200020025699200140001A15000017F0051D0F837324E00",
INIT_0B => X"5514554485D000000124002400000000000001004010A8812831605DA0000A05",
INIT_0C => X"708E2CB5320018CAC99BA0A3B9320018CAAAADA0C343F1AC1B01040A00202489",
INIT_0D => X"E7A3EE59320018CAC99BA0ACB9320018CAAAADA0CC421CA003B694B68018FAAA",
INIT_0E => X"24352AB2449A3FF2FA04E5E09B128834ADB1443A1891E4A928C29020E6A8524C",
INIT_0F => X"714C902375B801324301AB0067622E5E5404B2A5A40B1E6644AF0F021EA003AC",
INIT_10 => X"1216F50A8C241815FEB6A9158863F638FB60ED838E890B703C6260D8E3A21275",
INIT_11 => X"555E4C15F11133D171727A2550EE2F1BA0064F70DBDB1C74424E91E1C194C71D",
INIT_12 => X"ACCC59432A2B2D001F803471A9A960E57245FDF9D364DBD9435A6D45C9E81BED",
INIT_13 => X"0012CAC00006B0800000038814B72AB01508150013F162119014204373517700",
INIT_14 => X"002912300208092B940192D1000000000000A8A5AA80018120E0006600000000",
INIT_15 => X"1100011000110001100011000108000880008000520228080108039501200848",
INIT_16 => X"012000081500008A422150884081AC9000010003561180063DB4F61100011000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"28A28A3D2DE5F87963445469E79E7853D44C690DA64C1C69818768A360400000",
INIT_1B => X"F4FA3D3E8F4FA3D3E9A29A29A29A29A29A29A29A29A29A29A29A29A28A28A28A",
INIT_1C => X"000FA7D3E9F4FA7D1E8F47A3D1E8F47A3D1E8F4FA7D3E9F4FA7D3E9F4FA7D3E8",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"43FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE005500000000000000000000",
INIT_1F => X"80020005D2A95410FFFFC00000804154AA5D00001EFF78428AAA007BC2145F78",
INIT_20 => X"AD157400007BEAAAAAAAE955555D5568A105D2E974BAF7FBEAB45FFFFC00BAF7",
INIT_21 => X"007FC2000F78000010552E800AA002E821FFA2AAAAA00000417555FFD17DF45A",
INIT_22 => X"A08043FEBA5D55575FFF7AABFE00557BD74AAAAD17DF45F7D1421EF0055400AA",
INIT_23 => X"10FFD56AAAA5D043FFFFAAAABDEAA557BFDE00FFD140155F7AABDF55F7AE820A",
INIT_24 => X"FEF08517DF55A2FBEAB555D04154BAA2FBE8B55FFFFD55FF557FC2000FF80154",
INIT_25 => X"0000000000000000000000000000000000000000007FFDF45FF84000BA552ABD",
INIT_26 => X"28A821C7BC516DFF8438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE1049000",
INIT_27 => X"BE8B55FFF1C70BAF78A000005D2097438FFF1C7038140012482550E021C7EB80",
INIT_28 => X"0E1757DEBD17FF6DAADB504001C71EDA82AAA0955455D556DA00492490492F7F",
INIT_29 => X"3DF471C70851400BA0071C5028FF84020285D2085092002A801FFB6AAA8A1008",
INIT_2A => X"EBA4BAF6DE3AA8709208043FEBA555B555FFE3AABFE005D71D5492BED17FF45E",
INIT_2B => X"7557BC0028E38412428EBD16DA82410A3FFD7AAA4B8E824971F8E38E3DF45155",
INIT_2C => X"7DEB8000092552ABFFEF08517DF6DB6FBE8B555D04124BAB6FBE8B45E3FBD55D",
INIT_2D => X"55555003DE000000000000000000000000000000000000000000000000071FFF",
INIT_2E => X"00105D2A80145AA842AA00557BD75EFF78428B55AAD168B55F7FFFDFEFFFAA95",
INIT_2F => X"7FE10000000010F7FBEAB45FFD1554AAFFAE820105500154AAF7D5554BA55040",
INIT_30 => X"E801EFF7AEA8A10002E955FFA2D17DFFFAAFFC200055557DE00A280155455555",
INIT_31 => X"5557410F7D57DF55AAFBD55450055420BA0055574BAF784000BA5D0017410082",
INIT_32 => X"85568ABAA2FBD7545AA802ABEFA2AA9541000003DEBA557BD75EFA2AEBDE105D",
INIT_33 => X"FFFBEAB45AAFFD55555D7FC20AAA280000AAAAD17FE00082EBDF45AA8428A100",
INIT_34 => X"000000000000557FFEFA28402010552ABDFFF08517FFFFF7FBEAB455D04020AA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000002000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"5295B6957FCBE0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"6DE90201BF90102103AF158E805428249851BFB2C106592088DBF8400A5055C2",
INIT_05 => X"3824BD7F80148D9E07100A8201ED01C1A19B68F40A807ED9C18114956FF081DB",
INIT_06 => X"ED08CA6A8F033DD800000000050716BE9F57F8AC000807DFD999E0E5E1818B1B",
INIT_07 => X"00150886481240FE05A109228E2C0891D772A6F40045B8CF30E085DD2ED57D4E",
INIT_08 => X"72637FDF23800005981C0338190549C904182B6113870022000488C08B46268A",
INIT_09 => X"3E7437823DF78CDB6CA60E0E28EFFE2061872F80C1684A80C8604085F0074D3B",
INIT_0A => X"F5B4FFBD2FAD7FE653C36A1FF33E0E001E000B3A5DAADAFDDA5DA79350CFB801",
INIT_0B => X"CFE833C5C3D00018006C681700000000000000020012E9E10A31EB5FF9296A67",
INIT_0C => X"0D5ECE542A6FEEB2533EA160782A6FEEB2333EA16031F2BD47BDA2CA5D8164FC",
INIT_0D => X"282400F82A6FEEB2533EA160782A6FEEB2333EA160391BEFF2C32FB695F91911",
INIT_0E => X"573FAD5A86840354D1706FFFA3EF6E24B6D18C0D06638A207CFDE1F7DDAD76D5",
INIT_0F => X"FE4ACA4D77FAAB77CE3AF3EE78F58DB737E6E43E59AFE4A59B57679D19EFF2C7",
INIT_10 => X"ADB55572CA52606DFED6CA55334C04C04FF7D7A0ABD6DAAAB96529382B74E4E1",
INIT_11 => X"F9956EAA1A184045D5D7A870D2F5A5D7522D1281017F056E9C9C3FC95949C157",
INIT_12 => X"1F432EA58949D5B5C85F97871876F7D7E859FDEB974F486905001FDF5FA0D719",
INIT_13 => X"DEF20670021EE341036BF368128419FB5560158015177F916A039EF41FDB34A9",
INIT_14 => X"00633F1D0A7CC9AE7A08BFF0001D35682AC0CE8FCCC200A59BDD2FFE3F3EC7C7",
INIT_15 => X"FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A7800617112E46F05D02DD814102F8",
INIT_16 => X"05F08000179C16DECF67F08BC02F9086000D9E8A3F06ABD73DBCF4FBCF4FBCF4",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"34D34D48C4986868DC800181D75D7445F009EDCC4052E92E0204114F981800C0",
INIT_1B => X"1A8D468341A8D46834D35D74D34D35D74D35D74D34D35D74D35D74D34D34D34D",
INIT_1C => X"0008D46A351A8D46A351A8D46A351A8D46A351A0D068341A0D068341A0D06834",
INIT_1D => X"0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"43FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF5500000000000000000000",
INIT_1F => X"8028A00F7843FEBA55043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE00550",
INIT_20 => X"804154AA5D00001EFF78428AAA007BC2145F7D568B45000002010552EBDF45A2",
INIT_21 => X"5D2A95410FFAE800105D2A95410002A95410AAAEBFF55AAFFC00BAF7FFC00000",
INIT_22 => X"FFFD57DE00F7AE800AAAAAABDFEF5D2E974BAF7FBEAB45FFFFC00BAF78002000",
INIT_23 => X"AA5D517DF45AAD157400007BEAAAAAAAE955555D5568A105D7FFFFEFA2D568BF",
INIT_24 => X"1FFA2AAAAA00000417555FF8028B55082A974105D003FF55F7802AAAAAAD168A",
INIT_25 => X"0000000000000000000000000000000000000000000000010552E800AA002E82",
INIT_26 => X"955C71C043FE10490A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD749000",
INIT_27 => X"E050384124BFF7DB68A28A38F7803DE82490438FC7E3F1EAB55B6DF6DBFFF7AA",
INIT_28 => X"F5C70BAFFF1C7038140012482550E021C7EB8028A821C7BC516DFFDF68B551C0",
INIT_29 => X"FF1C70BAF78A000005D2097438FFAA85000492495428082E95400AAA0BDF7DB6",
INIT_2A => X"497FFAFFFB6D56FBFFEBDB78E38F7AA800BAB6AEBDFD75D2490492F7FBE8B55F",
INIT_2B => X"DEB8028AAAB6D16FA8249517FF6DAADB504001C71EDA82AAA0955455D556DA00",
INIT_2C => X"285D2085092002A801FFB6AAA8A10080E1757DEB8A2DB5514249243841003FF6",
INIT_2D => X"0BAF7FFFDF550000000000000000000000000000000000000000000000004020",
INIT_2E => X"8B55F7FFFDFEFFFAA9555555003DE00002ABFFEFF7FBFDFFFAAD168B55AA8000",
INIT_2F => X"D75EFF7FBEAB45552E954BA08003DFFFFFAAA8AAAF7843FE10000428B55AAD16",
INIT_30 => X"E95410AA843FFFFF7D5554BAF7D5554BA5504000105D2A80145AA842AA00557B",
INIT_31 => X"0000010F7FBEAB45FFD1554AAFFAE820105500154AAF7AE974000800154AA002",
INIT_32 => X"2801554555557FE10007FEABEFFFD57FFEFAAFFE8ABAFFAA820BAF7AEBFF5555",
INIT_33 => X"5500020AA08003DFFFA28028AAAF7D17DE0000517DFFFAAFFC200055557DE00A",
INIT_34 => X"00000000000004000BA5D0017410082E801EFF7AEA8A10002E955FFA2AABFF45",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000067FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"080BA868803F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"42016B0C401F58495C900A4859552A611D9A640F5903B2388004004C08A06008",
INIT_05 => X"16226B107811422A641C08038040007060E0032801E0202000991B708280B501",
INIT_06 => X"120886B3B8E0FC86142B4142B0000000011114D3058240240907F82000000000",
INIT_07 => X"006880802102401015610A02C4005000EA019D002482043FCF1C8090C02800C0",
INIT_08 => X"11018020D40A5004003260F9810541494D403D9B98810A0002C601000054B94A",
INIT_09 => X"022E0C6070000504102805C820C8016C30C250080C0182183804012A0A102200",
INIT_0A => X"084001E000108010230495A800FD865421432121804021C20452880C2D100000",
INIT_0B => X"3F140FC2060014250B9080008306C18360C1B0609C05013065CC042004040808",
INIT_0C => X"DF7C728582081483ACC15F9C3982081483CCC15F9CBA45505640000A40201900",
INIT_0D => X"DFEBFBF982081483ACC15F9F3982081483CCC15F9FB1962FCB69E08AAAEAEBCD",
INIT_0E => X"CAA02FE3F8E7F5E3AC3620805298B15A3FEBF1CFFF7670ACC3811A28AB57523C",
INIT_0F => X"01BD67DC4041D4CF03138DD865103EFEEAC9002BF05800D875E63CC9962FCB52",
INIT_10 => X"0016EA8DB7BFE25208E8F46A228BF8A757F1B72A8A800B7546DB9F1CA320037F",
INIT_11 => X"81A8A29509EAAE7FD3B749471C48F8A45981CCFAFDBF9464006FD037AEFAE515",
INIT_12 => X"EFF5778802A3AF8E8FB0440CE78773B709641256EC844B8AF92FD7CEDC24A9E1",
INIT_13 => X"0003C1C284601C2864000080113307E4800297D086E00036D2440E0880AAD62B",
INIT_14 => X"C44C92A88DCC2211E44174112840880000060D7030C30B885200D27400400808",
INIT_15 => X"0030800308003080030800308001840018400400602A01880980037109700C04",
INIT_16 => X"6808348340000020301805002D008CD943626111C0D95C20C2030A0030800308",
INIT_17 => X"C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B0",
INIT_18 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06",
INIT_19 => X"00000000000000000041B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_1A => X"1451451223059150A2EFB05C104104B3CEB80EE173C2300FCA8B7DF160000000",
INIT_1B => X"4AA552A954A25128955545145145155555545145145155555545145145145145",
INIT_1C => X"00025128944A25128944A25128944A25128944A25128944A25128944A2512894",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"43FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA0000000000000000000000",
INIT_1F => X"8400145AA801741000043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF550",
INIT_20 => X"7FBE8B45AAD568BFFFFAA975FF00003FE0055043FFFFFFFFFDFEFA2D56AB45AA",
INIT_21 => X"F7843FEBA55557FFEFA2D168B55AAFBFFFFFFF80021EF0855421EF00043FFFFF",
INIT_22 => X"A5D2A82155F7AEBFEBAFFD56AA00A2D568B45000002010552EBDF45A28028A00",
INIT_23 => X"BAA2FFC00000804154AA5D00001EFF78428AAA007BC2145F7D5400000004020A",
INIT_24 => X"410AAAEBFF55AAFFC00BAF7AE80010082E954BA0004174AAAA8428B45082ABFE",
INIT_25 => X"0000000000000000000000000000000000000000002E800105D2A95410002A95",
INIT_26 => X"00038F7DB6FBD7490E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA55041549214000",
INIT_27 => X"1F8FD7AAD16FB6DBE8E00155BE8015410140A3FFFFFFFFFDFEFE3F5FAF45AA80",
INIT_28 => X"5B471C7140438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE1049043FFEFE3F",
INIT_29 => X"124BFF7DB68A28A38F7803DE82495B78FC7AAD56FB6DBEF1FAFD7E384001EF14",
INIT_2A => X"FFD1420381C0A02082492A85155E3A4BDE92FFD56FA28B6DF68B551C0E050384",
INIT_2B => X"ABE8E28B7D1420BDEAAA2F1C7038140012482550E021C7EB8028A821C7BC516D",
INIT_2C => X"00492495428082E95400AAA0BDF7DB6F5C70BAFFAE870280024904BA1400174A",
INIT_2D => X"4BA550415410550000000000000000000000000000000000000000000002A850",
INIT_2E => X"DFFFAAD168B55AA80000BAF7FFFDF55002ABFFFFFFFFFFFEFF7FBFDFFFF7AA97",
INIT_2F => X"3DE0000043DFEFA2D56AB45AAD57DFEFF7AA82155F78015400552ABFFEFF7FBF",
INIT_30 => X"568B55A280021EF557FD7555550428B55AAD168B55F7FFFDFEFFFAA955555500",
INIT_31 => X"FBEAB45552E954BA08003DFFFFFAAA8AAAF7843FE10007FEAB55A2D17FFEFFFD",
INIT_32 => X"A842AA00557BD75EFF7D1400AA5D2A82000002A95545A2843FE00F7D17FEAAF7",
INIT_33 => X"0004020AA5D04154BAF7AEA8BEF55003DEAAA2D5554BA5504000105D2A80145A",
INIT_34 => X"0000000000002E974000800154AA002E95410AA843FFFFF7D5554BAF7AE974BA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000002000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000010228001000000000000000000024001620280000000000354200004008",
INIT_04 => X"00016200001310090090004840004152C7208802590000388000004C08006000",
INIT_05 => X"1621008008100002641C0803804000702000000000E02000009900000000B100",
INIT_06 => X"00A0010210200C00000000000000000000000080000000000000D82000000000",
INIT_07 => X"010084C00D267001B880080700285020020AC988200228024004804050089011",
INIT_08 => X"0E0E00000000000000106009872048400C4000010D000008000204150A00815A",
INIT_09 => X"022A040000000000000004C80000002C30C20000000002180800580000000000",
INIT_0A => X"0007600000000000000000080025860000000080A00020602040800000000000",
INIT_0B => X"031400C002000000000000000000000000000000000000000000000000000084",
INIT_0C => X"28DC0D385598035D0008A003B05598035D0008A0034078104B41A41000000000",
INIT_0D => X"041124505598035D0008A000B05598035D0008A0004263C0343EDD4140040422",
INIT_0E => X"B740500401180DE053A98F6ECC739D8140040231068187C39F5A4F985C008902",
INIT_0F => X"000010227848D4303807FC8CC5508AEAED1BFBD406451B02000E033263C0343C",
INIT_10 => X"D6480000000018A700FCF980CC300318A2420851546B2400000040D8549B5800",
INIT_11 => X"81C21140E40511802208D6B30C48F8A8A452210402120A936B0000000004C2A8",
INIT_12 => X"F9E9410006362A2B6424287B08286208D6B1427ED430B41402D0250823597001",
INIT_13 => X"0002C040000000000000000010030060009C000018440021011821B35254E99A",
INIT_14 => X"000040002000044000000000000000000002F0001F00002024B2000200000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"00000000000000000000000000008C8000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C30C30D0A208C4DC822EC1534D34C01FA3F0C7010C6600A0200441920000000",
INIT_1B => X"26130984C26130984C30C30C30D34C30C30C30C30D34C30C30C30C30C30C30C3",
INIT_1C => X"000130984C26130984C26130984C26130984C26130984C26130984C261309A4D",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D00000000000000000000",
INIT_1F => X"AA974BA5D517FFFF08043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA007",
INIT_20 => X"FFFFFFFFF7FBFDF55A28402000F7D56ABFF557BFFFFFFFFFFFFFFFFFBFDFEFFF",
INIT_21 => X"AA8017410007BFFFFFFFFFFFFEFF7D16AB45AA8002000F7D5575455D043FFFFF",
INIT_22 => X"5AAD568B55F7AE955FFAA840201008043FFFFFFFFFDFEFA2D56AB45AA8400145",
INIT_23 => X"FF5D043FFFFF7FBE8B45AAD568BFFFFAA975FF00003FE00557BFFFFFFFFBFDF4",
INIT_24 => X"FFFFF80021EF0855421EF002ABFFEFF7D168B55AAD17FFEFF7AE975FF00557FF",
INIT_25 => X"000000000000000000000000000000000000000000557FFEFA2D168B55AAFBFF",
INIT_26 => X"954AA5504154921471FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA55000008255000",
INIT_27 => X"FFFFEFF7FBFAFD7E3A4954BA555B7AFC7080E3FFFFFFFFFFFFFFFFBFDFEFFFAE",
INIT_28 => X"DF52545550A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD74975FFFFFFFF",
INIT_29 => X"AD16FB6DBE8E00155BE8015410147FFFFFFF7FBF8FC7EBD568B55A28000000FF",
INIT_2A => X"497BFDFC7E3F1FAF55A2DB6FB7DF7AE955C7BE800000008043FFEFE3F1F8FD7A",
INIT_2B => X"7EBA0955FF145B7AFC7410438FC7E3F1EAB55B6DF6DBFFF7AA955C71C043FE10",
INIT_2C => X"C7AAD56FB6DBEF1FAFD7E384001EF145B471C71424B8FC7E3D56AB6DB6DF7AFC",
INIT_2D => X"4AA550002000550000000000000000000000000000000000000000000005B78F",
INIT_2E => X"FFEFF7FBFDFFFF7AA974BA55041541055517FFFFFFFFFFFFFFFFFFFFEFF7AA97",
INIT_2F => X"FDF5500517FFFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB45002ABFFFFFFFFF",
INIT_30 => X"56AB55A28002000F7FFC2155552ABFFEFF7FBFDFFFAAD168B55AA80000BAF7FF",
INIT_31 => X"043DFEFA2D56AB45AAD57DFEFF7AA82155F78015400557BFDFEFF7FBEAB55A2D",
INIT_32 => X"FAA9555555003DE00007FFDF45AAD568B45AAFBFFFFFFFAA95545F7840201000",
INIT_33 => X"AAD16ABFFFFFBEAB45A280155EF557FE8B55000428B55AAD168B55F7FFFDFEFF",
INIT_34 => X"0000000000007FEAB55A2D17FFEFFFD568B55A280021EF557FD755555042AB55",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000004000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"0001E6000053300B00D0005800000000000000407B0004BB830004DC3D01E000",
INIT_05 => X"FEE0000008720043EC3C3D0F87FA19F7E0201C409BE1F10623BB000A100CF300",
INIT_06 => X"00200006102FFC8E0007C00078008000171175A200096404D97FFBE4744200AA",
INIT_07 => X"000000482491301000010001DC00000000000000004203FE4005800000008030",
INIT_08 => X"40800020E2008000027FEFF946058180010429000001080AAA010F8000000000",
INIT_09 => X"03EAFE400000120000913FD80000003DF7DE0080010047FBF8000000000800C5",
INIT_0A => X"0800000080000010000400080FFDBE0000004000000100000100506002204610",
INIT_0B => X"FF14FFC00600000000801020000000000000010240001721214E000004000000",
INIT_0C => X"A70C0008020000200000000F30020000200000000F3008001E00000000001803",
INIT_0D => X"004A58F0020000200000000F30020000200000000F3040200000020000000026",
INIT_0E => X"000000000019B140000800800000020000000030B86000400080000200000000",
INIT_0F => X"000014AC08000000508001030A0A4001000000000002183E61E6000040200001",
INIT_10 => X"0000000000A56000090100000000001F86C00010080000000000525801000000",
INIT_11 => X"0600000000001716800000803102020000000002BC360020000000000292C010",
INIT_12 => X"06049CDF70C08040100000706707600000801000000000000057450000100106",
INIT_13 => X"000ADFC011001C81080001101F977FE008000000000000400400400020000805",
INIT_14 => X"0000000000000000000000020020029000000000000000020000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000002000200000000",
INIT_16 => X"0080800801810100000000000093ED8000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000401",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"18618640C49821201C0001A1E79E79A4B0038200010089054C1A0104D2040020",
INIT_1B => X"0C86432190C86432196596596596596596596596596596596596596586186186",
INIT_1C => X"00086432190C86432190C86432190C86432190C86432190C86432190C8643219",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA5504020100800000000000000000000",
INIT_1F => X"AA974AA550002000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7",
INIT_20 => X"FFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFFFFFFFFFFFFF7",
INIT_21 => X"5D517FFFF087FFFFFFFFFFFFFFFFFFFFDFEFFFAE974AA5D003FE005D043FFFFF",
INIT_22 => X"FF7FBFDFFFAA84000105D556AB55557BFFFFFFFFFFFFFFFFFBFDFEFFFAA974BA",
INIT_23 => X"EF08043FFFFFFFFFFFFFF7FBFDF55A28402000F7D56ABFF55003FFFFFFFFFFFF",
INIT_24 => X"B45AA8002000F7D5575455D2EBFFFFFFFFFFFEFF7FBEAB55A28000010F7D16AB",
INIT_25 => X"0000000000000000000000000000000000000000007BFFFFFFFFFFFFEFF7D16A",
INIT_26 => X"954BA550000082557FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA55040002800000",
INIT_27 => X"FFFFFFFFFFFDFEFF7AE974BA5500050380071FFFFFFFFFFFFFFFFFFFFFFFF7AA",
INIT_28 => X"0038E285D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA55041549214043FFFFFFF",
INIT_29 => X"7FBFAFD7E3A4954BA555B7AFC70871FFFFFFFFFFFFFFF7FBFDFFFFFAA974BA55",
INIT_2A => X"490E3FFFFFFFFFDFEFF7F1FAFC7A28002028555F6FB7D5D75FFFFFFFFFFFFEFF",
INIT_2B => X"5A28402010FFDB6ABEF140A3FFFFFFFFFDFEFE3F5FAF45AA8000038F7DB6FBD7",
INIT_2C => X"FFF7FBF8FC7EBD568B55A28000000FFDF525455524BFFFFFFFBFDFC7E3F5E8B4",
INIT_2D => X"4AA5504000BA080000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFEFF7AA974AA550002000557FFFFFFFFFFFFFFFFFFFFFFFFFFAE95",
INIT_2F => X"1541055043FFFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08517FFFFFFFFF",
INIT_30 => X"FFFFEFF7AE974AA550028AAA5D2ABFFFFFFFFFFFEFF7FBFDFFFF7AA974BA5504",
INIT_31 => X"517FFFFFFFBFDFEFFFFFEAB45AA80154AA557BEAB4500557FFFFFFFFFDFEFF7F",
INIT_32 => X"A80000BAF7FFFDF55002EBFFFFF7FBFDFEFFFD568B55A284020BA557FFFFFF5D",
INIT_33 => X"F7FBFFF55A2D16AB45AA8402000F7FBEABEF5D2ABFFEFF7FBFDFFFAAD168B55A",
INIT_34 => X"0000000000007BFDFEFF7FBEAB55A2D56AB55A28002000F7FFC215555043DFEF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"1094EC681244819000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"0001E6000053300F01D4587800446194F49020107F0012BBC00202DC3823EA82",
INIT_05 => X"FFF201B228704123FC3C381F87C03DFFF012412A9FE1E01013BF09404050F300",
INIT_06 => X"100B3096F43FFF002004020044041084CB01AD0000037617027FFFE050000080",
INIT_07 => X"A12034043C802A821D41412001A0040950AB60014114C3FE4187A009A663A680",
INIT_08 => X"7F40002C01004000047EFFF811A46968004060629A0002208A00000068113205",
INIT_09 => X"E3EBFE0A812D8D5B742D3FF84056383FF7DE0880042107BFF9C45B85101C49A3",
INIT_0A => X"02804A08221890004806C0310FFDFE00040009814C089202225412115414601D",
INIT_0B => X"FF56FFC0281280080180B2948004400220011100841200D001000624000100C0",
INIT_0C => X"50025360694101816002D41A4068C101815004D8158809C86065941840B1014F",
INIT_0D => X"82418A0068C101816002D41A40694101815004D815810D42E04A08A80098C024",
INIT_0E => X"1A300012682960828F05C96A001B029010134160C8125B0B271802242880A044",
INIT_0F => X"49F115100920C54E8EA256ECF078BA081C10080E05C0B06AA8B12CFD0D42E044",
INIT_10 => X"5144104F30A8801406D00290006280320100010362A8A20826A88660D86B2020",
INIT_11 => X"8010602011819E290048A2118EC8140C08064802C0081B0D64040936443306C5",
INIT_12 => X"C322A4C40A0300600C0A80509F418008804581BA0038005A706680012280506A",
INIT_13 => X"18DBFFC000120080002341881F3FFFF80DCC158092C044600466208CC5091011",
INIT_14 => X"806520398C6021569249C4B3007127080806FF917FC30010107688862A28C545",
INIT_15 => X"9228D9228D9228D9228D9228D99146C9146C84006309044081A001B188300E20",
INIT_16 => X"0448008004000000E07008010003EF80022A51904595123203040D9228D9228D",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_19 => X"0000000000000000004010040100401004010040100401004010040100401004",
INIT_1A => X"7DF7DF7FEFFDFDFFFBE7F3FCF3CF3FFF6EFF7FFDF7FF3EFC1FBFFDF7E0000000",
INIT_1B => X"FEFF7FBFDFEFF7FBFDF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF",
INIT_1C => X"001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFD",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D00020000800000000000000000000",
INIT_1F => X"AE954AA5D00020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"55000200000003FFFFFFFFFFFFFFFFFFFFFFF7AA974BA5D0402000557BFFFFFF",
INIT_22 => X"FFFFFFFFEFF7AE974BA5D00174BA00003FFFFFFFFFFFFFFFFFFFFFFF7AA974AA",
INIT_23 => X"BA5D043FFFFFFFFFFFFFFFFFFFFEFF7AE954BA5D04174AA00003FFFFFFFFFFFF",
INIT_24 => X"FEFFFAE974AA5D003FE005D2EBFFFFFFFFFFFFFFFFFFDFEFF7AE954AA5500174",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFD",
INIT_26 => X"974AA550400028007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000001000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"04050005571FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082557BFFFFFFFF",
INIT_29 => X"FFFFDFEFF7AE974BA55000503800003FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5D",
INIT_2A => X"140E3FFFFFFFFFFFFFFFFFFDFEFF7AE954BA5D00154AA00043FFFFFFFFFFFFFF",
INIT_2B => X"FFFAA974BA5D00104925D0E3FFFFFFFFFFFFFFFFBFDFEFFFAE954AA550415492",
INIT_2C => X"FFFFFFFFFFFF7FBFDFFFFFAA974BA550038E285D2ABFFFFFFFFFFFFFFFFBFDFE",
INIT_2D => X"4BA5D00000100000000000000000000000000000000000000000000000071FFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02000557BFFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7FFFFFFFFFFF",
INIT_30 => X"BFDFEFF7AE954AA5D041740055517FFFFFFFFFFFFFFFFFFFFEFF7AA974AA5500",
INIT_31 => X"043FFFFFFFFFFFFFF7FBFDFEFFFAE954BA5500174AA08043FFFFFFFFFFFFFFFF",
INIT_32 => X"7AA974BA550415410552ABFFFFFFFFFFFFFF7FBFDFFFFFAA974AA5D00174BA08",
INIT_33 => X"FFFFFDFEFF7FBFFFFFF7AE954BA5D0000010552ABFFFFFFFFFFFEFF7FBFDFFFF",
INIT_34 => X"000000000000557FFFFFFFFFDFEFF7FFFFFEFF7AE974AA550028AAA5D2EBFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"8632CA211E4491D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"24B000808800040439245B221373581F97B0A8D1040F92000F42000047A00E58",
INIT_05 => X"011B2BBA308F023810004700083E220811E9BF2844021B1004045E4249500449",
INIT_06 => X"EF018980A51003AA0200C020088E16A85235722940A817251100040D6D0702A2",
INIT_07 => X"24E8145C9ECAB0D247B013B405EAD525FAE48FC2060B880081A26DCD4047EFF9",
INIT_08 => X"0050482D0141C0055280100751096B6A40D6F86723E510AA2004803D3275EB20",
INIT_09 => X"20110204804818CD280100207246A8020000AC0283002004051507A5411C0DA0",
INIT_0A => X"4E506A2C6898B2950AA6D635B00041C23020131A80CFDFF3FE509A907C556828",
INIT_0B => X"002200050F60E220A06880D2A14050A028501428054278142151262CA5034385",
INIT_0C => X"F06273612B3482C0C0078E1F412B1582C090078E1F840A2B0114020104022460",
INIT_0D => X"C2C0DB012B1582C0C0078E1F412B3482C090078E1F891C239F8908003099C1AC",
INIT_0E => X"0828041BA859F213AFC14AA380430060181BA1B0FD16770236A4091621C08055",
INIT_0F => X"095337B08AA600CA88B143AB11880C280600101F09C030AB28B03C111C239F87",
INIT_10 => X"3096004B61BD8068B92400D0004E30368910E8822A984B0025B0DE6089462660",
INIT_11 => X"F07830001AC2173B00E162563454C40804055412D4481128C4CC012A66F30455",
INIT_12 => X"BF006850840180A00E1C81900C4190E160589C48082C006A9057CA4385809520",
INIT_13 => X"39C020004416B105036B4180C000800C8C00460848952220592745AC11A544B1",
INIT_14 => X"103D2A512C6A8C4F0008AA800470370000A0004D0000002126F30C902A29C545",
INIT_15 => X"C2A81C2A81C2A81C2A81C2A81C9540E1540E001400006100003202D040050220",
INIT_16 => X"45E22022365034A8EA754008004C0214202C50013456520CA09281C2A81C2A81",
INIT_17 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_18 => X"0040100401004010040100401004010040100401004411044110441104411044",
INIT_19 => X"0000000003FFFFFFFF9004010040100401004010040100401004010040100401",
INIT_1A => X"3CF3CF7FE7FDFD7DF7EFFDDDF7DF7DF7DEFE8FF1F7DEBD6FCD9F7DF7D0512289",
INIT_1B => X"FE7F3F9FCFE7F3F9FCF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"0007F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04000000000000000000000000000",
INIT_1F => X"AE974BA550000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D00020AA5D7FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D00000AA007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAA954BA5504000AA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA",
INIT_23 => X"BA5D7BFFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500020BA5D7FFFFFFFFFFFFFF",
INIT_24 => X"FFFF7AA974BA5D040200055517FFFFFFFFFFFFFFFFFFFFFFFFAA954BA5500000",
INIT_25 => X"000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040200008000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"00020BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAA954BA5D00000BA557FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5D",
INIT_2A => X"5571FFFFFFFFFFFFFFFFFFFFFFFFFAA954BA5504020AA5D7BFFFFFFFFFFFFFFF",
INIT_2B => X"FF7AA974AA5D00070925D71FFFFFFFFFFFFFFFFFFFFFFFF7AA954BA550000082",
INIT_2C => X"FFFFFFFFFFFFFFFFFFEFF7AA974AA5D040500055517FFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D040200008000000000000000000000000000000000000000000000003FF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAA954AA5D00020AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA5504",
INIT_31 => X"7BFFFFFFFFFFFFFFFFFFFFFFFF7AA954BA5D00000BA5D7BFFFFFFFFFFFFFFFFF",
INIT_32 => X"7AA974AA55000200055517FFFFFFFFFFFFFFFFFFFFEFF7AA974BA5504020BA55",
INIT_33 => X"FFFFFFFFFFFFFFDFEFF7AE974AA5D00154105D517FFFFFFFFFFFFFFFFFFFFEFF",
INIT_34 => X"000000000000043FFFFFFFFFFFFFFFFBFDFEFF7AE954AA5D041740055557FFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"5886C0201A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"0005EE040057700F40D08078500000D9218020407F0000BB8018A2FC380BEAC2",
INIT_05 => X"FFE0419028700023FCBC385F87C0BFFFE0124002FFE1E0C517FF09111212F300",
INIT_06 => X"DF0AF116D03FFC96102081020000020489019C4304802412027FFFE000000000",
INIT_07 => X"B710000001160A003475C8100123400E20E1F40F439647FF4807E189A477EF81",
INIT_08 => X"7F0F94801008000007FEFFFB110140695812CC4188D58A0AAA10803448D0844F",
INIT_09 => X"C3EBFD4201258112D4487FF8001010FFF7DE4000000003BFF8C2581808002001",
INIT_0A => X"0801000C024000004A9400000FFDFF50010103134CAFDF03BA18000F39900037",
INIT_0B => X"FF57FFC02812F00429DC92C40002000100008000105400C00400100000A01800",
INIT_0C => X"424202A1CAF13F214001521001CBF03F21100152100801C17E61841950B1C10F",
INIT_0D => X"420B8001CBF03F214001521001CAF13F2110015210088528E00E02C8200A430A",
INIT_0E => X"12480202C86040902AC60BACDF0E02D02001C1C044006D0C94FB94320880603C",
INIT_0F => X"09B00300010AF5052419D196441902801430182800A018D9CA8000648528E00D",
INIT_10 => X"C140004D101808458A5602E000892029110445C19960A00026880C0067390000",
INIT_11 => X"4040301009408021144CB042F880100C0601844068880CE72000013600600332",
INIT_12 => X"EE38A1F80E02120018390320F050144CB241D0B9023402085020825132C8CB5B",
INIT_13 => X"001BFFC200400020224000405F7FFFE0008E17C0D240406519400500840A9524",
INIT_14 => X"907120AC810033149249C433200180082A06FF907FC308181204800600000000",
INIT_15 => X"1010C1010C1010C1010C1010C10086080860840063090442A18001B188300C48",
INIT_16 => X"2000100100000000000004002403EFC10302219A41C1443243050C1010C1010C",
INIT_17 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_18 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_19 => X"0000000000000000000080200802008020080200802008020080200802008020",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"550000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974AA550400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"00087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550402010087FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE954AA5D00000AA007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA5504020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974AA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA55",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400010087FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE954AA5D0402038007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550400028",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE954AA5D00020BA087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"00010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA550002010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D00",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974AA550002000087FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE954AA5504000BA087FFFFFFFFFFFFFFFFFFFFFFFFFFAE954AA55040001000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAA954AA5D04000AA087FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007BFFFFFFFFFFFFFFFFFFFFFFFFFAA954AA5D00020AA007BFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"0000745C200801000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"0001E6000053300F00D0007810042140C00000407F0000BB800000DC3801EA00",
INIT_05 => X"FFE0000008700003FC3C380F87C019FFE01240009BE1E00003BF00000000F300",
INIT_06 => X"DC8C3006103FFC0000000000000000048900880100800012027FFFE000000000",
INIT_07 => X"0061200009B24B043980021000810284204A8001401643FE4007E5501AA00000",
INIT_08 => X"7F00000000000000007EFFFB11A56940581280031D61420000B080102040BC5B",
INIT_09 => X"C3EBFC020125811254083FF80000003FF7DE0000000003BFF800580000000001",
INIT_0A => X"0580000000000000000000000FFDFF4000000AA0354000019C40000128000011",
INIT_0B => X"FF56FFC000104000000010440000000000000000001000C00000000000000240",
INIT_0C => X"48C0804012500021B00880108012500021E00880104809C1666594584031010F",
INIT_0D => X"0501840012500021B00880108012500021E0088010492064206100E810842000",
INIT_0E => X"0270040410004C840041A0D8005410903804100144800803419043064900C002",
INIT_0F => X"400041020902F60002260D65B361BAA1041018140F02C0000809408D20642053",
INIT_10 => X"D0021800020818B06D9802F00030C02060110002C9E8010C00010480B35A0300",
INIT_11 => X"90203020042108603100061516EE800C060228204300166B4060080008240593",
INIT_12 => X"14AE4C7C02000040206602C10B48110006143B62023C00142800B04400095DFF",
INIT_13 => X"001BFFC000000000000000001F17FFE000DC1180C78044000440292083010402",
INIT_14 => X"814080008000010012414433000100080806FD107FC300000000000600000000",
INIT_15 => X"1000C1000C1000C1000C1000C100060800608400630104408180012188300C00",
INIT_16 => X"0000000000000000000000000003EF80020201904181003003000C1000C1000C",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"3DF3DF64C7986120B42BB99575D75FFD2AF6E7CC1132CD73DF3A441990000000",
INIT_1B => X"1E0F0783C1E0F0783DF7DF7DF7CF3CF3CF3CF3CF3DF7DF7DF7DF7DF7DF3DF3DF",
INIT_1C => X"0000F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100800000000000000000000",
INIT_1F => X"AE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"00007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0002000087FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D00020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0400010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA550002000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0000010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA550002000007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010080000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0000010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D000001008",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA550000010087FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA550002010087FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00004000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"4909E6093253306F82D0007C80000000080E01007F8020BBC00040DC3801EA00",
INIT_05 => X"FFE0000008704503FE3C380F87C019FFF01241009BE1E00203BF80800000F392",
INIT_06 => X"CC083006103FFF9E2086C2086E006604C9019D03108B7412027FFFE070400880",
INIT_07 => X"0000004024057000000100000000000000000001401643FE4007C00000000000",
INIT_08 => X"7F00000801404000007EFFFF40010000401408000045000000A0801000408000",
INIT_09 => X"C3EBFF4A7DF795965C6D3FFC0020003FF7DF01880C618FBFFDD75E0010004043",
INIT_0A => X"0000000000000000009400000FFDFFC006020000000000019804000028000191",
INIT_0B => X"FF56FFC02812E0182000F2C48304418220C11160845004D04820000000000000",
INIT_0C => X"0800800002400001000800000002400001000800000801C0786184185031810F",
INIT_0D => X"0400000002400001000800000002400001000800000000202000000800000000",
INIT_0E => X"0200000000000404000000880000001000000001000000000090000008000000",
INIT_0F => X"000040000100C600800001040000040009100000000200200000400000202000",
INIT_10 => X"4000000002000000081001000000000040010000082000000001000001080000",
INIT_11 => X"0000400080000040010000001080001008000000010000210000000008000010",
INIT_12 => X"0420000000030280000000010000010000001020000000000000100400000108",
INIT_13 => X"001BFFE0120012C1400080291F17FFF0018C11808200400000400000C2000000",
INIT_14 => X"80400000800001001243443B000100880806FD107FC301800000000600000000",
INIT_15 => X"1000C1000C1000C1000C1000C10006080060840077330C4889CC292588300C00",
INIT_16 => X"44C82082068C0200000008014023EF80020201904189003003000C1000C1000C",
INIT_17 => X"4110441104411044110441104411044110441104411044110441104411044510",
INIT_18 => X"1104411044110441104411044110441104411044110441104411044110441104",
INIT_19 => X"2FFFFFFFFFFFFFFFFFC110441104411044110441104411044110441104411044",
INIT_1A => X"0924821409005312E8A25E15A69A6BFB0A196A8C5A2932F7C13C15DA08080000",
INIT_1B => X"C46231188C462311892492492492492492492492482082082082082082092482",
INIT_1C => X"00162B158AC562B158AC562B158AC562B158AC562B158AC562B158AC562B1188",
INIT_1D => X"0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"00087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04000",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0400000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402000",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040200000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402000087FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0400000007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"94A7B2B1450000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"6FEBEF5FEC737AFBC6F85FDEB220109E1FEFFFE3FBA7FDFB9BD301DC3FF5F0D2",
INIT_05 => X"FEEDBFDC387F987FEF7C3FAF87FF59F7F5FB7FF59BE1FF980BBBB7FE6D21F3DB",
INIT_06 => X"DFA08957902FFDEE9D7DC9D7DF2B263893479DDFAFDFE15213FFFBE1F1D3A333",
INIT_07 => X"00018010992310605CE10301DE0C1831CB7DF60A244B9BFEE00589DDBCEFEDC1",
INIT_08 => X"FFEFAA001D8EA111DA7FEFF90F21C8C84D9C0D858FC7020828C18FD18346BBF0",
INIT_09 => X"0BFAFFF37DF7B9DF7DCB3FDE89ECC07DF7DF5F985C6BCFFBFA28F99E7EB07F47",
INIT_0A => X"0607307DCFE1D4077B4D0026FFFFBE7D67D7F3BB79CFFB83BF14EC1E7D598058",
INIT_0B => X"FFFCFFC7D7D51D6F5FDCB935D7AFEBD7F5EBFBF7FEBD66DBFCA3F87501AE7B08",
INIT_0C => X"40520201F45EC0010007E01001F45EC0010007E010084BCD7FF1B61B5C33813F",
INIT_0D => X"0001A001F45EC0010007E01001F45EC0010007E01001BD8020500008001F0100",
INIT_0E => X"0200001EC00040B02007EC09A0E00010001DC0004600400F781429C008000077",
INIT_0F => X"81C203404B3BFD0402346235408402C08010003C064000E408010081BD802060",
INIT_10 => X"68B1000E401A08FE0012040000FC002001360403E434588007200D00F88C84C0",
INIT_11 => X"281D00001F01002156040675809145400007B00040091F1190982038406807C8",
INIT_12 => X"903A80008320C0403C34000088601604067D00212000007C400082D81009FC08",
INIT_13 => X"D6BFDFF7BFFED3FBFF6A84383F177FF005FFBFF5FA1040076065F730FC08043A",
INIT_14 => X"CDEBCFF589807B7096CD4CF73AC1FC98884FFF19FFC71FEFED7B251E35768E8E",
INIT_15 => X"78C0D78C0D78C0D78C0D78C0D7A606BC606B8C56F7730ECCDBDF152199F51EDD",
INIT_16 => X"FEFDFDDFE7DD87FEFF7FF796FFFFFDFFD7E681B867D3683A03A40F78C0D78C0D",
INIT_17 => X"EBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFB",
INIT_18 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAF",
INIT_19 => X"6FFFFFFFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_1A => X"4C30C375E2BD54D5D6C565F871C71D44FCF491E166CC853E8695F86EDB5C8864",
INIT_1B => X"26130984C26130984C30C30C30C30C30C30C30C30C30C30C30C30C30C30D34D3",
INIT_1C => X"000130984C26130984C26130984C26130984C26130984C26130984C26130984C",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"1085B0B041000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"6FAB975B6470BAF386C87A9CB00000001FEF9F23E3A7BDE79B5101D23FB5C0C2",
INIT_05 => X"F8EDBFD4347F18778E723F2E47FE59C7F5FB7F759B91FB880BA3B6FE2921CBDB",
INIT_06 => X"DFC00147000FFC128D5CE8D5CC210638A046889CAB57E84217FFE3E181932377",
INIT_07 => X"000141000000042000000288020C18300320620A80231BFE200181092CE7ED80",
INIT_08 => X"FEEF22000C562551D87E8FF90041101042110180004102800008801183468180",
INIT_09 => X"0BE0FC137FF7A0FF75813F1C85244071EFBF17D85C738BE3FA08F9DE36B05B07",
INIT_0A => X"040510768EA0C406630D00226FFE3E2D62D6E21259CFDB039E806C0245188040",
INIT_0B => X"FF48FFCC57550D63564D1D2556ADAB56D5AB6AD7EAB962CBD8A3A83101F47E08",
INIT_0C => X"00130201E44A40010007600005E44A4001000760000843C561E5C55C42B9011F",
INIT_0D => X"00002005E44A40010007600005E44A40010007600004BD8020100008001F0100",
INIT_0E => X"0200001EC00000382006EC0820A00010001DC0000208400D781020C008000077",
INIT_0F => X"81C20040431BC50402146235400400408010003C064000C400018080BD802020",
INIT_10 => X"4821000E400204FE0010040000FC0000003E0403A424108007200102E8888080",
INIT_11 => X"080500001F0100005E040475808101400007B00000015D111010203840081748",
INIT_12 => X"903A8000012040403C34000080201E04047D00202000007C400000F81001FC08",
INIT_13 => X"109E1FE5ADA4C25ADE72041A3F147FF0018DBBB5FA10400360649310FC08003A",
INIT_14 => X"EFABC7054880693016DD4C755AC16C1A884FFE18FFD757E7ED7A211E81C09818",
INIT_15 => X"3440C3440C3440C3440C3440C3C2061A2061AD46FF730E5CCBCD55219AB55F0D",
INIT_16 => X"DE75ED5EC71385FC2512E3565BBBF1BAD6F281BC63F1683803C00E3440C3440C",
INIT_17 => X"AB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6B",
INIT_18 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6AD",
INIT_19 => X"7FFFFFFFFFFFFFFFFFAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_1A => X"0000003C010072F24388521000000140A8100481CA8604368714104A47168874",
INIT_1B => X"8040201008040201000000000000000000000000000000000000000010400000",
INIT_1C => X"00140A05028140A05028140A05028140A05028140A05028140A05028140A0100",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201008",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010087FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"8C2100804900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"02000100440408002408008002221000204116A280000F000001400000100010",
INIT_05 => X"0004D44400004D4400000000000000000000005C0000000A0000002C20600000",
INIT_06 => X"2000004100000120040A0040A00B009000620294010000400080000888800911",
INIT_07 => X"2488045002489020420110800244891211440804000810002000081040000000",
INIT_08 => X"00B062080542C004CA00000050080202008401842004108AAAA00008912240A1",
INIT_09 => X"2800010000000C0000E400002040500000009202C10020400044000222000204",
INIT_0A => X"02043058C460540329810002D002000400407020800000004000640800088008",
INIT_0B => X"0008000140000401028008330000800040002002480102010082981500062108",
INIT_0C => X"00500000040A40000000A00000040A40000000A0000040060084104110828030",
INIT_0D => X"00012000040A40000000A00000040A40000000A0000000800010000000000000",
INIT_0E => X"00000000000000A00000040020A000000000000006000000080020C000000000",
INIT_0F => X"8000024040152000000020000004004080000000000000240000000000800020",
INIT_10 => X"0821000000120002000004000000000001220000040410800000090000808080",
INIT_11 => X"0805000000000001420000200001014000000000000900101010200000480008",
INIT_12 => X"0000000001204000000000000820020000200000200000000000028800002000",
INIT_13 => X"29400000933050080C0001900020000000408010000000022000D61028000008",
INIT_14 => X"440245400082D022040000400800081022C0000080000206CB0821082B694D4D",
INIT_15 => X"605016050160501605016050160280B0280B0012000843066021001400040024",
INIT_16 => X"0810840861CD33548542A10209D4100E4040A00002002C004001036050160501",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008021",
INIT_18 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_19 => X"0000000000000000000020080200802008020080200802008020080200802008",
INIT_1A => X"41041001A835050788440B58C30C31DF6C110A00246972C0C39989A40A0C22E1",
INIT_1B => X"C06030180C060301810410410410410410410410410410410410410410410410",
INIT_1C => X"00160B0582C160B0582C160B0582C160B0582C160B0582C160B0582C160B0180",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"00000000000000000000000000000000000007FFFFFFFF800000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0803B2814D0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"26E1E905CC574828C4F85FC600000016004F77E2F887CDB80BC340DC07D1F000",
INIT_05 => X"FE1DFE4C080F884FE33C078F803F19F011E93ED49BE01F1A03B8972E6D20F049",
INIT_06 => X"64A08857902000DE142D4142D5030010134395D70589415002FFF800F0C38111",
INIT_07 => X"00088400092300601CE00101DE040811D919F402244293FEE00400CCB46BA4C1",
INIT_08 => X"7FA0AA08148A4000887FE0000F20C8C80D080D818FC2000000418FD08142BAD0",
INIT_09 => X"0BFA02E204D2154D28AA3FC60888D03C10415A80402847F8002458926A002E45",
INIT_0A => X"0406305587A1540231410006DFFF80540541619968C76980E914E4163D498010",
INIT_0B => X"FFFC0007C7C0140D0B50A8218102C0816040B1225C1506512C83E85500AC3A08",
INIT_0C => X"40520000141EC0000000A01000141EC0000000A01008480D3EB4A24A0C910037",
INIT_0D => X"0001A000141EC0000000A01000141EC0000000A0100100800050000000000000",
INIT_0E => X"00000000000040B000010401A0E000000000000046000002080429C000000000",
INIT_0F => X"80000340483B590000202000008402C080000000000000240801000100800060",
INIT_10 => X"28B10000001A08020002040000000020013600004414588000000D00108484C0",
INIT_11 => X"281D000000000021560002200011454000000000400902109098200000680088",
INIT_12 => X"000000008320C00000000000086016000220000120000000000082D800082000",
INIT_13 => X"D6ABC032936E43A92F2880B01F37001004B29450580000066021F6303C000408",
INIT_14 => X"45624DB481806A62840800C22800B8900042FF0180000ABFEF89250815568A8A",
INIT_15 => X"68D0068D0068D0068D0068D006A68034680300021410028450530014014002D4",
INIT_16 => X"2C989489418D13FE7F3FFD8BADB7FC4F4164A00806522C0A40A50268D0068D00",
INIT_17 => X"C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C4B1",
INIT_18 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02",
INIT_19 => X"2FFFFFFFFFFFFFFFFFC0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_1A => X"5D75D7FFEFFDF9FAF3E7E3EFFFFFFEBFD6EE7FFDF7FE78FC3CEFFDFFEA0C0060",
INIT_1B => X"EFF7FBFDFEFF7FBFDF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DD75D75D7",
INIT_1C => X"001F7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDF",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"3CF3CF75EFBD75F5FFEFFDFDF7DF7FFFFEFF9FE1F7FFBFEFDFBBFDFFD0000000",
INIT_1B => X"FE7F3F9FCFE7F3F9FCF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"0007F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"1084B030000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"6DA986092050306382C05A1C900000001FAE89016387B2A38B5000D03FA1C0C2",
INIT_05 => X"F8F92B90307F41338E303F0E07FE19C7F1FB7F289B81FB8003A396D20940C3DB",
INIT_06 => X"DF800106000FFC020004C0004C0006288004880800036002137FE3E101030222",
INIT_07 => X"000100000000000000000220000810200220620E00030BFE000181092CE7ED80",
INIT_08 => X"7E4F400000000001107E8FF90001000040100000004102200000801102448100",
INIT_09 => X"23E0FC027DF780DF74013F1C00240071E79F05888C618BA3F800599C10104903",
INIT_0A => X"040100240A808004420400202FFC3E002202021259CFDB039E00080245100000",
INIT_0B => X"FF40FFC407500020004C10060204010200810040801060C04821202001A05A00",
INIT_0C => X"00020201E04000010007400001E0400001000740000803C0616184184031010F",
INIT_0D => X"00000001E04000010007400001E04000010007400000BD0020000008001F0100",
INIT_0E => X"0200001EC00000102006E80800000010001DC0000000400D7010000008000077",
INIT_0F => X"01C200000308C50402144235400000000010003C064000C000010080BD002000",
INIT_10 => X"4000000E400000FC0010000000FC000000140403A020000007200000E8080000",
INIT_11 => X"000000001F01000014040455808000000007B00000001D010000003840000740",
INIT_12 => X"903A8000000000403C34000080001404045D00200000007C400000501001DC08",
INIT_13 => X"001A1FE004048240426200081F147FF0018C1380DA10400140640100D4080032",
INIT_14 => X"812982050800A91012494C31004124080886FE187FC301B124F2001600000000",
INIT_15 => X"1000C1000C1000C1000C1000C18006080060840477330C4889CC012188310E08",
INIT_16 => X"44602002061004A820104809402BE1900222019861D1403803800C1000C1000C",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"2FFFFFFFFFFFFFFFFF8100401004010040100401004010040100401004010040",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000100080",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000007C01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000",
INIT_1E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020100000000000000000000000",
INIT_1F => X"AE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007",
INIT_20 => X"FFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_21 => X"5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFF",
INIT_22 => X"FFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA",
INIT_23 => X"10007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFF",
INIT_24 => X"FFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04020",
INIT_25 => X"0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF",
INIT_26 => X"974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000000",
INIT_27 => X"FFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE",
INIT_28 => X"0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFF",
INIT_29 => X"FFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D",
INIT_2A => X"007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFF",
INIT_2B => X"FFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010",
INIT_2C => X"FFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFF",
INIT_2D => X"4BA5D0402010000000000000000000000000000000000000000000000007FFFF",
INIT_2E => X"FFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE97",
INIT_2F => X"02010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFF",
INIT_30 => X"FFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D04",
INIT_31 => X"7FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFF",
INIT_32 => X"FAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D040201000",
INIT_33 => X"FFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_34 => X"0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFAE974BA5D0402010007FFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


end;