library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_master is
	port(clk             : in  std_logic;
        address_a       : in  std_logic_vector(31 downto 2);
        enable_a        : in  std_logic;
        wbe_a           : in  std_logic_vector(3 downto 0);
        data_write_a    : in  std_logic_vector(31 downto 0);
        data_read_a     : out std_logic_vector(31 downto 0);

        address_b       : in  std_logic_vector(31 downto 2);
        enable_b        : in  std_logic;
        wbe_b           : in  std_logic_vector(3 downto 0);
        data_write_b    : in  std_logic_vector(31 downto 0);
        data_read_b     : out std_logic_vector(31 downto 0));
end; --entity ram     

architecture ram_master of ram_master is
signal enable_a_lo       : std_logic;
signal wbe_a_lo          : std_logic_vector(3 downto 0);
signal data_write_a_lo   : std_logic_vector(31 downto 0);
signal data_read_a_lo    : std_logic_vector(31 downto 0);
signal enable_b_lo       : std_logic;
signal wbe_b_lo          : std_logic_vector(3 downto 0);
signal data_read_b_lo    : std_logic_vector(31 downto 0);
signal enable_a_hi       : std_logic;
signal wbe_a_hi          : std_logic_vector(3 downto 0);
signal data_read_a_hi   : std_logic_vector(31 downto 0);
signal enable_b_hi       : std_logic;
signal wbe_b_hi          : std_logic_vector(3 downto 0);
signal data_read_b_hi    : std_logic_vector(31 downto 0);
signal address_a_reg     : std_logic_vector(31 downto 2);
signal address_b_reg     : std_logic_vector(31 downto 2);
signal enable_a_lo_256       : std_logic;
signal wbe_a_lo_256          : std_logic_vector(3 downto 0);
signal data_write_a_lo_256   : std_logic_vector(31 downto 0);
signal data_read_a_lo_256    : std_logic_vector(31 downto 0);
signal enable_b_lo_256       : std_logic;
signal wbe_b_lo_256          : std_logic_vector(3 downto 0);
signal data_read_b_lo_256    : std_logic_vector(31 downto 0);
signal enable_a_hi_256       : std_logic;
signal wbe_a_hi_256          : std_logic_vector(3 downto 0);
signal data_read_a_hi_256   : std_logic_vector(31 downto 0);
signal enable_b_hi_256       : std_logic;
signal wbe_b_hi_256          : std_logic_vector(3 downto 0);
signal data_read_b_hi_256    : std_logic_vector(31 downto 0);
begin
process(clk)
begin
if rising_edge(clk) then
	address_a_reg <= address_a;
	address_b_reg <= address_b;
	end if;
end process;
data_read_a <= data_read_a_lo when (address_a_reg < x"0001000"&"00") else
data_read_a_hi when ((address_a_reg >= x"0001000"&"00") and (address_a_reg < x"0002000"&"00")) else 
data_read_a_lo_256 when ((address_a_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_a_hi_256 when ((address_a_reg >= x"0003000"&"00") and (address_a_reg < x"0004000"&"00"));
data_read_b <= data_read_b_lo when (address_b_reg < x"0001000"&"00") else
data_read_b_hi when ((address_b_reg >= x"0001000"&"00") and (address_b_reg < x"0002000"&"00")) else
data_read_b_lo_256 when ((address_b_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_b_hi_256 when ((address_b_reg >= x"0003000"&"00") and (address_b_reg< x"0004000"&"00"));
enable_a_lo <= enable_a when (address_a < x"0001000"&"00") else '0';
enable_b_lo <= enable_b when (address_b < x"0001000"&"00") else '0';
enable_a_hi <= enable_a when ((address_a >= x"0001000"&"00") and (address_a < x"0002000"&"00")) else '0';
enable_b_hi <= enable_b when ((address_b >= x"0001000"&"00") and (address_b < x"0002000"&"00")) else '0';
enable_a_lo_256 <= enable_a when ((address_a >= x"0002000"&"00") and (address_a < x"0003000"&"00")) else '0';
enable_b_lo_256 <= enable_b when ((address_b >= x"0002000"&"00") and (address_b < x"0003000"&"00")) else '0';
enable_a_hi_256 <= enable_a when ((address_a >= x"0003000"&"00") and (address_a < x"0004000"&"00")) else '0';
enable_b_hi_256 <= enable_b when ((address_b >= x"0003000"&"00") and (address_b < x"0004000"&"00")) else '0';
wbe_a_lo <= wbe_a when  enable_a_lo='1' else x"0";
wbe_a_hi <= wbe_a when  enable_a_hi='1' else x"0";
wbe_b_lo <= wbe_b when  enable_b_lo='1' else x"0";
wbe_b_hi <= wbe_b when  enable_b_hi='1' else x"0";
wbe_a_lo_256 <= wbe_a when  enable_a_lo_256='1' else x"0";
wbe_a_hi_256 <= wbe_a when  enable_a_hi_256='1' else x"0";
wbe_b_lo_256 <= wbe_b when  enable_b_lo_256='1' else x"0";
wbe_b_hi_256 <= wbe_b when  enable_b_hi_256='1' else x"0";



ram_bit_0_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"441406267B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"0005802424830120024121209088809DF81454ACA01E03501D0A3B91E00F0A00",
INIT_05 => X"E0F001CC00012034C20B0232838F80D001C0100AEC83C008EF101A034C8CC300",
INIT_06 => X"2F1620F1721BA346AA2C95C5CB1400000161F84322000DA8C40F003C80030780",
INIT_07 => X"5939F36677EE1C387777622717EF711004A6818111086008E080FDC305940018",
INIT_08 => X"13160400195E83A3A0F61BC3929ECB622AABF5FF83860CEB164833F179B48CEE",
INIT_09 => X"01036D8004FDB47600000229410C61010016DC998C84B0128202C0DCB48F05D5",
INIT_0A => X"4400402A0A37000182502440888420247041E876810099D35F900002DB00105C",
INIT_0B => X"AD4434020CA2E0B32B01A752B078412A24818094151348062400E2A034D86444",
INIT_0C => X"3E2781EA781E2781EA781E2781EA781E2781C33C0613C0E21028840239452116",
INIT_0D => X"394818429A95E954868AD0E52273F54258000080808900C3807122C3E04E0338",
INIT_0E => X"8E3B15C94001120055704DC4A1624487E2489024481224091282C4300942A194",
INIT_0F => X"C06101C55D65C3E3F01F52FFC1E0013C1F801F52FFC1E0013C1F8090423D38A1",
INIT_10 => X"ECC381C0118796BE001F567FC1E0013C1F801F567FC1E0013C1F9085DFBF7E15",
INIT_11 => X"F885DFBF7E30F00C0270F3751F1FD00FECBF7E25C0700463E17B2C7F811FD7AD",
INIT_12 => X"C40FE6474190626D6491063597F9177B956EF378D33E4030061341F077C571F8",
INIT_13 => X"0C4DAE207F328E3082636B2807FFD80FE00007E03F7207D3E03F9167184131B5",
INIT_14 => X"1F4FE047EFA0CAE06101C53E3647D3F144FCDD22B81C0098E57D9081FCE8C852",
INIT_15 => X"38574FF31ADF08DBF81846A540049707E0FE3307D3F141FFB45478040570EED4",
INIT_16 => X"90240902C189601208A1102B4AA5584B4068000019A80098120BCA4C617635C9",
INIT_17 => X"0240902409024090240902409024090240902409024090240902409024090240",
INIT_18 => X"2409024090240902409024090240902409024090240902409024090240902409",
INIT_19 => X"9AA09426A8000000000000000009024090240902409024090240902409024090",
INIT_1A => X"104104104104431042720EE38E38AAF9A93E7131C136AD8E9B562CF03B2E8E78",
INIT_1B => X"F87C3E1F0F87C3E1F0F87C104104104104104104104104104104104104104104",
INIT_1C => X"FFC00001F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0",
INIT_1D => X"AAAAABDEBAF7AE8000000000000000000000000000000000000000000000C200",
INIT_1E => X"EFF7D142145A2AE800BA08514214555517DEAA5D7BFFEAAF7803FEBAF7FFD74B",
INIT_1F => X"E00A2FBD75FFFF84001550851555FF55517FE000055421FF00557DF45A2D5401",
INIT_20 => X"74BA552EBDFFF0004020005D5555555A2AABFFFF5D516AA00A28028A00AAAEBF",
INIT_21 => X"3FEBA082ABFE10AAAEA8ABA55517FF45A2AEBDEBAAAAAA8BFFF7D140010FF841",
INIT_22 => X"FD75FF0051401FF5D00154105504000BA5D2E97545A28028B450855401450804",
INIT_23 => X"FBFFF45A2FFFDE00002E801FFA2AABFE00FFFFD74AA085540000002E801FF557",
INIT_24 => X"0000000000002ABEFAA80001EFF7FFC20BAF7D1575450800020BA08517FF45F7",
INIT_25 => X"57803AEBAF7F5D74AAA2A03AA38BF8FC00000000000000000000000000000000",
INIT_26 => X"7A3F00516DA2D5451D7EBDB47155BC2A87092AAFA9257F1C5BC00AA5D7FF8EAA",
INIT_27 => X"00EA8000150A801C01C7142EBFBC7EB8005B55A85B555EF095F50578085BE8FC",
INIT_28 => X"BEAE3D542A004380124921D20975FFAAA1521FF492BF8F40B6AAB84AF555168A",
INIT_29 => X"8F6DE05B40480557A95A3A1C2EBAE28168ABAA2D43D568BC5400168E90E2F412",
INIT_2A => X"47B50A80095178157FEFA0742FA3AA28EA8168A954100071D2E90A855C7A00A3",
INIT_2B => X"0A8F57F6DA971F8F7FFFA42D16D1EAE925EA0BFEBF4AA09217F4905684170851",
INIT_2C => X"000000000000000000000000000002D57AAA8402A8743DBD202DA95568A95E80",
INIT_2D => X"17D34ABA5D7BEAAAAD786BCEAAFFD1564BA2282BFA02A2C28000000000000000",
INIT_2E => X"007F8B2B2D97D483AFA7BD9F5EFA87F57555AAFBD7555FFAE95408A8FDC31AD0",
INIT_2F => X"0A6AEA8FAF0451CA001D4845C2087383F79A5046A37B55F38415555797D63BFF",
INIT_30 => X"A7D7463CC508D07577BAFBD542000D382964A92B401E71D7581C33172EC0A030",
INIT_31 => X"0502828811FCD4EABDB1DFDFC8365A2FD5E04AA5780A8AAAD7AC3CA02003BEBB",
INIT_32 => X"4FF72AAADF245595157050790621F562B1122DA70C3808458881056A5502AA15",
INIT_33 => X"F6A03D4BFB79AFA4C5CB5F5896D55BBAAC55EAFAF86D35E4A92B4460D1506037",
INIT_34 => X"FC0000007FC0000007FC0000007FC0000007FC0000007FC07AAF12E00505D3FD",
INIT_35 => X"7FC0000007FC0000007FC0000007FC0000007FC0000007FC0000007FC0000007",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000400000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"650C00000848A0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000004208B00200E010800006667BE7000102C00080000040012010000080C",
INIT_05 => X"0080000000002020600100208D04414000800000000200004800080000800200",
INIT_06 => X"04022140220932C2038900000100000008082010000000800488000000020400",
INIT_07 => X"088C0060242183060CF118011281B00000220010400020002081A00082100001",
INIT_08 => X"40000400014812466427040098C000622AAAA43E3060C158AC97F0356BDBFBD0",
INIT_09 => X"00026C000559102400200281400469000008B0800000901080004004308B4340",
INIT_0A => X"045413002200000000400408200000201041000208000040020820034200005C",
INIT_0B => X"41E11C008089540000420100101088400000808404004000000020A000100414",
INIT_0C => X"18C191AC191A4191A4191AC191AC191A4191A00C8560C8D08400000609010100",
INIT_0D => X"0E08A20BC417C16004C0B8382210904018000080100100012200000064064019",
INIT_0E => X"0E0615C96000000010200000802100022008100408020401020040100142200E",
INIT_0F => X"C06100000021E300B000000781E00140018000000781E00140018000002430E3",
INIT_10 => X"68C381C00000024E0000000781E00140018000000781E0014001908400005E11",
INIT_11 => X"088400003C30F00C000000155800D00000003E21C0700000000F001180000004",
INIT_12 => X"4000260640900004A400081401A0000004041218503E40300600000048043180",
INIT_13 => X"00009A0001208C30800025200003D807E0000000007252016000904618400013",
INIT_14 => X"480160000F00C0E06100000012D2005100409520381C00000005920004C0C812",
INIT_15 => X"0004025000120850B8180625400400000010711200510004B414780400000055",
INIT_16 => X"1004010040002002080000000804000A0000000011A000100208C008611430A0",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"5800050008000000000000000001004010040100401004010040100401004010",
INIT_1A => X"1451451451564090C69606492492C09A8C205148D757DF8A94102E0001063A29",
INIT_1B => X"BADD6EB75BADD6EB75BADD555555555555555555555555555555555555555145",
INIT_1C => X"FFE0000174BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974",
INIT_1D => X"F5D2AAAB555555400000000000000000000000000000000000000000000303FF",
INIT_1E => X"EFA2D17DEBAF7D1574BAAAFBFDFFFA2FFD74000855555FFFFFFC01FF087BE8BF",
INIT_1F => X"145557BFDEAA5500154AAAAAEBFF455D04175FF5D7FEAAAA002ABDEAA5D2EBFF",
INIT_20 => X"20BAAAD540145F7D5574BAAA8415400005540155F7D16AB45002EA8ABA005540",
INIT_21 => X"975EFF7AEBFF550055555FF55003DE00A2FFFFFEFAAD57DE00082AAAA00082A8",
INIT_22 => X"16AABAAAAEBFE10AAFBD7545F7D5554AA5D2ABDEBA082A821455D2EA8B455D2A",
INIT_23 => X"FFEABEFA2FBEAB455D7BD55FFFF84155FFFFFFFFF55AAAABFFFF5D556AB45A2D",
INIT_24 => X"000000000000175FFF7D140010FF84174BA552EBDEBA0004020AA5D04155FFAA",
INIT_25 => X"4BFBC51FF1471E8BEF55242FF47015A800000000000000000000000000000000",
INIT_26 => X"0B6AEBAEAA5D2EBDFFFBED17FEAAF7D5524AAA2F0BAF7FABDFC7E10005F525D7",
INIT_27 => X"55142A8708202FBD257F1C7550492490E17EAAA2AAB8F4515043DFC75575C700",
INIT_28 => X"03D1420AD000B420820AAE2DB6FB6DF7DFD5038ABA140A2D00554517DEBDB6FB",
INIT_29 => X"25555F8FFDE38087FC51C7F7AABFF55BC5B555C74B8A38E38085BE8B47A3A005",
INIT_2A => X"BA4AF555168B68FEDF6AB52AAABD21EF1C2FEA5FDEBDB505FA4920AFE10082E9",
INIT_2B => X"17AEB8BFF155552B6F5E8BFF1EFBFDBFF5FF1C00BF5D25475C7B7FEAFF45BEAA",
INIT_2C => X"00000000000000000000000000000151EAE3D542A004380124921D20BFFFA0AA",
INIT_2D => X"3D795000087BC01458AFBC11FF55516ABEFDD003EFE5093DC000000000000000",
INIT_2E => X"550434D555C53E0CE2AAA8742BA5D2ABDFFFF7D57DEAAFFD5420B2A2D37DB07A",
INIT_2F => X"F0851575FFAAFBDD5542B2EDD608897FD610D01151C610592A974BAFBAC28B55",
INIT_30 => X"100F3D68FFFAABAC20EF04003FE102400144ABAAFFF7DE772FDD56588042F72E",
INIT_31 => X"4EA0006BFE007E2E8315DD02F6A81A239501755F504BDF557D79431FD006EABA",
INIT_32 => X"03158517BD745AEAEA8FAF0C55EAF57FF957CAAA7FABF7DFD0C6A7DFFFA07FC0",
INIT_33 => X"964A92B403EE18D5408A6F2AFADF6900FFFF68BEFDFFB4B1FE5551141E78A028",
INIT_34 => X"0000000000000000000000000000000000000000000000165BAFBD542000D382",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000400000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0812",
INIT_01 => X"2145A00A1079284D04A044A54E504368404000720885800802000006ECD10200",
INIT_02 => X"5C010800020408040C415854AA055254090541A111000A104A00000009083510",
INIT_03 => X"0C1000100C0000D40526480250149120031500A0218808002440804288890550",
INIT_04 => X"8840C28120051400582012021808040409C0B26850488419444010C10A024A49",
INIT_05 => X"488510910548012025C0C0000300086854B141042252142042A048D090006372",
INIT_06 => X"948037480159A403109848000428AA8282102040449090D520085224410AA420",
INIT_07 => X"01020402242000408468112010810C055200022025A83AA3008882004A001542",
INIT_08 => X"11491C154429220A2824640010A010020282843E0008124C0000211000008840",
INIT_09 => X"E280442C1411D020828A2B116824632885419240016001900AE01A2020066395",
INIT_0A => X"30105108880684145002021012D40D718241108815380200900160AE42CE2818",
INIT_0B => X"53419F10308D100054AA080092112C100B400880454058E80B94080C49318000",
INIT_0C => X"D0090D0090D2890D0890D2890D0890D2090D0048610486808403A384880B8981",
INIT_0D => X"8202043800000620500403080A919000B8AD0304144008111A00582043243050",
INIT_0E => X"9835300002AA40AA902408200010002021060C810241832241280C81A0984020",
INIT_0F => X"100000000080A0000140000002000140200A8000000200014020100290E469C6",
INIT_10 => X"00100000000003400A8000000200014020094000000200014020087000000000",
INIT_11 => X"014200000004000000000081400004C00000000020000000008C000010A00000",
INIT_12 => X"0510000000000006800001880004008400800000000020000000000048100000",
INIT_13 => X"0000D0260000000000003409280000000000000040025000030000000000001A",
INIT_14 => X"400002A0000000000000000042900000A100000000000000008012A200000000",
INIT_15 => X"000000004420300000000000000000000010C010000098000000000000000105",
INIT_16 => X"00802208036408C0820010004D36A222120090554000E40080000000088000A0",
INIT_17 => X"8802008020080200822088220882208802008020080200822088220882208802",
INIT_18 => X"8320883200812008120081208832088320883200812008120082208822088220",
INIT_19 => X"E88051029FC0FC0FC1F81F81F820883208832088320081200812008120883208",
INIT_1A => X"08208208208C13A4301040B2CB2CBAC838B6C0080271AE180616A851158E2863",
INIT_1B => X"944A25128944A25128944A082082082082082082082082082082082082082082",
INIT_1C => X"FFE381F928944A25128944A25128944A25128944A25128944A25128944A25128",
INIT_1D => X"A550002000AA800000000000000000000000000000000000000000000003C200",
INIT_1E => X"BAFFAE801FF087BE8BFF5D7BEAA1055042AA105555421EFFFD568AAA002EBFEB",
INIT_1F => X"FFFA2D57DE10557BE8ABAF7AAA8BEFAAAE975FFA2D5555450851574000851554",
INIT_20 => X"5555F7D568ABAF7D5574BA552EA8AAA5D2EBFFFFA2D1554BAF7D17FEBAAAFFFD",
INIT_21 => X"EAAAA552AAAAAAAAAABFF455D04175FFFFD5574AAAAAA974BA082EA8BEFAAD55",
INIT_22 => X"FEAA000055401555D7BFFE10085557410F7AA97410087BD55FF087FEAA10A2FF",
INIT_23 => X"0017400550402155A2803FE005D7FE8B45F7FBFDE00085540155F7D56AA00007",
INIT_24 => X"00000000000017400082AAAA00082A820BAAAD540145F7D557410AA8428A1055",
INIT_25 => X"4BD16FAAA002ABFEAA550E82000E28A800000000000000000000000000000000",
INIT_26 => X"FEAFBD2410005F57482E3AA801FF1471E8BEF5574AFA00010ABFA38555F401D7",
INIT_27 => X"AAF7D5524AAA2F1FAF7FABFBFF400417FEF082F7AAA8BEFE2AA955EFA2DB5757",
INIT_28 => X"492082EADBFFBEDB55555E3DF6DA82F7DF520385D2FE80AA5D2EBDFD7BED1574",
INIT_29 => X"21C7005B6FB47F7A438E925D24ADAAAB6AAB8F455784155C75575C7000B6AE95",
INIT_2A => X"4717DEBDB6FA3D0075EDA800051C05571474024A81C5557578EBA087400007FC",
INIT_2B => X"FFDE381D716FA15550015428E10A001FFB40038F68F7F578F7FFEF568E280855",
INIT_2C => X"000000000000000000000000000001043D1420AD000B420820AAE2DB4716DF7D",
INIT_2D => X"828FDEBA5D7BC015582D57DEAA002ABDEAA552A80010AAA88000000000000000",
INIT_2E => X"AAAE955EFAAFBC15F5A3D7D6800087BD5410AAAA801FF55556ABEF5D517EEE00",
INIT_2F => X"A5D2ABDF55F7D575EAAFFD50A2B2A3D169B07A3D7BFE10597BFDE00AEAC28BFF",
INIT_30 => X"555A53C00B2A2AA02000082ABDFEFFFFBC1154AAFFFFE107FF9D72A20842080B",
INIT_31 => X"4EAA28015400547FC315D00797CF4780286A2105D2A3FEBAFFAC28B555504145",
INIT_32 => X"99ADABD5A8AAA0051575FFA2FFFDA02003FFDEAA8557D65550915544AA5D5157",
INIT_33 => X"144ABAAFFD75E7F2BDDD2B8016F9E2555500174AA282E20BFFFF842AAAAADD56",
INIT_34 => X"0000000000000000000000000000000000000000000000030EF04003FE102400",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000800000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380206",
INIT_01 => X"200C9A40408001683C0462C99E004B61404040028804A0080A000416A0990A0C",
INIT_02 => X"4809A900031800444461089866E331352180D468B8040E600C0081110B802CD0",
INIT_03 => X"6D0B61108C00014231A3080408C68420330066010A80881068A808401CC46330",
INIT_04 => X"482218066A09C03B348C1C1928DD5A4402211A68470944842640902107002D24",
INIT_05 => X"0583180353202020000144E50B44644B30A86D05014A0D224063095092100E34",
INIT_06 => X"54023740216934020303680A040066D98A182210085A50C02048288234629414",
INIT_07 => X"018C00220430814204E01C581291820CCA000E3226413990008C80205A00CCCC",
INIT_08 => X"4108747320081246252D5010184000220002A43E10294258E805E1156002D940",
INIT_09 => X"D0AA546AC41B112029A61D84424429AA1320B1010140C1350B48292020024180",
INIT_0A => X"000102022850A1CC0047071913208CE802430488082042008040F399606F4058",
INIT_0B => X"5141BE42B88840005268081412152900484201A814144D60888CAA2C48151020",
INIT_0C => X"1B49019490194901B4901B4901949019C901B64805E480CA94480506980125C4",
INIT_0D => X"5A01E2B1080602E00C54216800859000199C98800C8140A11A44423040240450",
INIT_0E => X"28A65300E6664599902600009821204A040C1C040C0205038300480801480208",
INIT_0F => X"000000000090000003202900000010002008A02900000010002008039666928B",
INIT_10 => X"00000000000801000A202900000010002009E0290000001000200A3800008000",
INIT_11 => X"036000008000000000000088000002D003008000000000000280100016200812",
INIT_12 => X"05B008088000008201021C880000488002810005000000000000040000100000",
INIT_13 => X"0010402B80412000000410199800040000000000408020000680209000000208",
INIT_14 => X"800012980040300000000000C020000C8300208800000000008200AE01011000",
INIT_15 => X"40A0000841003100010401000000000002008020000C38000200000000000120",
INIT_16 => X"10070300704028820801400068360424820185CCE0128010020000008088021C",
INIT_17 => X"0070100701007010050180501805018050180501805018070100701007010070",
INIT_18 => X"070140601007014060100701C040180501C040180501C0401807010070100701",
INIT_19 => X"4A81454A26AA555AAB554AAB5541C040180501C040180501C040180501406010",
INIT_1A => X"08208208209441D0B0000092492480AA2860607818F18E0C851428200B262C31",
INIT_1B => X"D4EA753A9D4EA753A9D4EA492492492492492492492492492492492492492082",
INIT_1C => X"FFD55E21A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8",
INIT_1D => X"FAA8000155080000000000000000000000000000000000000000000000000200",
INIT_1E => X"EFFFD568AAA002EBFEBA555142000AA802AA10F7D57FEAA557BE8B45A2D5555E",
INIT_1F => X"A10550402000AAD56AAAA557BC0155A280021EFA2FFE8B4555042AA105555421",
INIT_20 => X"0010AA842AAAAFFD542000FFD5574000851554AAFFAE801FF087BC01FF5D7FEA",
INIT_21 => X"7DE105551420BAF7AAA8BEFAAAE975FF005540145A2D157410AAD17DFFF5D040",
INIT_22 => X"03DEBAAAFFFDFEFAAD57DEAAF7AE975FF080428B455D7FFDEAA5D55574BA0051",
INIT_23 => X"AE800AA087BD5555552A821EF007FFFEAAAAD5554AA552EBFFFFA2D5554BAF78",
INIT_24 => X"000000000000020BA082EA8BEFAAD555555F7D568ABAF7D5574BA552E800BAAA",
INIT_25 => X"E975EAB6DBEDF575FFAA8E02155080E800000000000000000000000000000000",
INIT_26 => X"5EBAEADA38555F451D7EBD16FAAA002ABFEAA555E02000E28AA8A38EBD578E82",
INIT_27 => X"FF1471E8BEF5575EFA00012A87A38AAD56DA824975C217DAA84021FFAAF5EAB5",
INIT_28 => X"400BED57FFD7410E05038BE8E2DABAFFDB47412ABFE90410005F57482E3AA801",
INIT_29 => X"FEBA5D71D742A407FFFE00555F47082E3AAA8BEFA02A955EFA2DB5757FEAFBD2",
INIT_2A => X"BFFD7BED157482F7803AEAAA2F1FAF7FABFBEAE2AEBA4974871C043AB6D4975F",
INIT_2B => X"F7AE38497FC00BAB6A4850821C75D25C74920821D708757AE2AA3FFC04AA552E",
INIT_2C => X"0000000000000000000000000000007092082EADBFFBEDB55555E3DF6DA82F7D",
INIT_2D => X"AA8A8ABAAAD568A1020516ABFFFFFFD75FFAAAE8014500288000000000000000",
INIT_2E => X"AA80001FFAAD57EB55A2A8ABEBA5D7BD5545A2D57DEAA002EBDEAA557BC0010A",
INIT_2F => X"0087BD5410AAAA801FF5555629EF5C517EEE00828D74AAFBD57DE000057C21FF",
INIT_30 => X"EFA8FBC15E5A3D5D7400FFD57DF55082E974AAFFAABDEBA77FDD66A0ABBDC200",
INIT_31 => X"50555002ABFF54517EEB25D57C14100957FF6105D7BD5400AAAC28BFFAAAE955",
INIT_32 => X"FA42A3D7020BA5D2ABDF55F7D1554A8FFC42AA10A7D169F57ABD7FEEBAAA8415",
INIT_33 => X"C1154AAFFFFE10FFF9DF202096F014AAFF84154105555C215500000014558557",
INIT_34 => X"000000000000000000000000000000000000000000000015400082ABDFEFFFFB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000400000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204002",
INIT_01 => X"01039802000820491C00650E1E004340403008418984014902030906A8D10200",
INIT_02 => X"480108A000000000444048E41E80F00A41043118680002000800000009882390",
INIT_03 => X"06504110080000D0040608024010102026001260300000003080880208C000F0",
INIT_04 => X"9100E98268154C1AE0B01C160033B944028290285AE0DC38E02090E81C22E801",
INIT_05 => X"5C0F20B36F000109200044C401041C4CF21C48B433483C8242EAE1B0000074C4",
INIT_06 => X"100007000059800310086A1A0022E18780000140C9D9D0930000F228075A6071",
INIT_07 => X"00000000242000008461000810818403C100060064012E00048C82201800BC28",
INIT_08 => X"0048CC8F01090602202C0400008000002202243E400010480000211540008810",
INIT_09 => X"40E0DC1EB5191120C7BE7D152201612E80E891E0614041340838450020422111",
INIT_0A => X"30545DAD8C2E0982400603003200872003FB1408082840002044007846164E0A",
INIT_0B => X"43411D10118D1A04522E000498140C104B260DA0404003C08B6000AC01128000",
INIT_0C => X"C5010C3010C1010C3010C1010C1010C3010C140869808618850BE6305989AB80",
INIT_0D => X"100140302800108018840440028480001B8780800000003102045C3443043410",
INIT_0E => X"3080620481E0E18790012A001001026808000002020101028100200180080201",
INIT_0F => X"000000000010000005C0200000001000000C4020000000100000000380E4C308",
INIT_10 => X"00000000000800000D00200000001000000EC020000000100000086A20008000",
INIT_11 => X"012820008000000000000008000001B00100000000000000020000002AA00010",
INIT_12 => X"06D0000080000080000241D80000800442800001000000000000040000000000",
INIT_13 => X"0010003A00002000000400021800040000000000008010000B00001000000200",
INIT_14 => X"400005900000100000000000801000089000008000000000000200F800001000",
INIT_15 => X"00000000A500100000000100000000000200001000002E000200000000000020",
INIT_16 => X"000000C032700000022400444934240A8021B63C005108010004100098098010",
INIT_17 => X"C010080200401008000040300800004010000200C01000020040100802004030",
INIT_18 => X"02000000000100C0300400008000000300C0100C00000020080000C030000000",
INIT_19 => X"20240142325930C9A6CB261934C000200801004030040200800000030040100C",
INIT_1A => X"14514514514E98264686668A28A260521CC45140C700FC0A0002870980831A28",
INIT_1B => X"1A8D46A351A8D46A351A8D555555555555555555555555555555555555555145",
INIT_1C => X"FFD5E7D8341A0D068341A0D068341A0D068341A0D068341A0D068341A0D06834",
INIT_1D => X"A5D55420AA002A80000000000000000000000000000000000000000000000200",
INIT_1E => X"AA557BE8B45A2D5555EFAAD140155080000155FF843FFEFAA84001FF5D043FEA",
INIT_1F => X"000AA80001555D04174AA002A80010FFAE975FFAA80001EFA2AAAAA10F7D57FE",
INIT_20 => X"00BA5D51555EF002AA8BFFAAAAAAA105555421EFFFD568AAA002EBFEBA555542",
INIT_21 => X"82000AAD568AAA557BC0155A280021EFA2FFE8B45F78400145FF842AAAAA2AA8",
INIT_22 => X"BC01FF5D7FEAA105D0428B4500003DFEF080428B455D002AABA5D2AAAAAA5D2E",
INIT_23 => X"80154BAA2FBE8AAAF7AA821EFAAAAA8BEF552E820000851554AAFFAA801FF087",
INIT_24 => X"00000000000015410AAD17DFFF5D0400010AA842AAAAFFD542000FFD57DF55A2",
INIT_25 => X"A284051D755003DE92415F42092142E000000000000000000000000000000000",
INIT_26 => X"71C0A28A38EBD57DE824975EAB6DBEDF575FFAADE02155080E85145E3803FFEF",
INIT_27 => X"AA002ABFEAA555F42000E2AA851455D0A124BA002080010FFA4955C7BE8E021C",
INIT_28 => X"145F7802AABAA2A480092415B505D71424AABD7F68E2FA38555F451D7EBD16FA",
INIT_29 => X"AA824924AAA92550A07038BED56DA824975C217DAA84021FFAAF5EAB55EBAE82",
INIT_2A => X"55482E3AA801FF1471C01EF5575EFA00012ABFB6D080A3AFEF080A2FB45490E2",
INIT_2B => X"B6FA12ABAEBDF7DAA80104BAAAFFEAA00F7AE821D7B6A02FBC71D0E10010005F",
INIT_2C => X"0000000000000000000000000000010400BED57FFD7410E05038BE8E2DABAFFD",
INIT_2D => X"02897555A2803FFFFAA841754555043FE10087BC2000552C8000000000000000",
INIT_2E => X"FF8017545F7AE821455D2CAAABAAAD57DE1000516ABFFFFFBD75FFAAFFC01450",
INIT_2F => X"A5D7BD5545A2D57DEAA002EBDEAA557BC0010AAA895555042E820BA080400010",
INIT_30 => X"FFAAD57EB55A2A880155F7802AAAAAA8002010007FC0155D5022A955FFACBFEB",
INIT_31 => X"BEF002EBDF45542AAAA0008043CAB0552C97CAAFFD57DE000057C21FFAA80001",
INIT_32 => X"CFE55D2CC2000087BD5410AAAA801FF5555421EF58517EAB00028A9BEF002EAA",
INIT_33 => X"974AAFFAABDEBAF7FDDE6A0AA90FDFEFA280020BAA2FFEAA10FFAE82145F7803",
INIT_34 => X"000000000000000000000000000000000000000000000002000FFD57DF55082E",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000800000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A337A20E07C0C1E006",
INIT_01 => X"295FBC468000A04D5C6A60000C34C24841280A00084000C8C212892EEAD53235",
INIT_02 => X"C809AD5CB118E640A4D158F8011FF0002080000082C8C66609DB7DDDCB1F2036",
INIT_03 => X"250906263A4C904214A35C80085285720B20648A88800000B8E0F852A884500E",
INIT_04 => X"4005122126899100064D20001044429C78A43A2C4436CC87198A3916E0551A24",
INIT_05 => X"A370C14CA0E900004048402389CFE2F20F7D7A354CB5C208E51437F044948912",
INIT_06 => X"9B9407B9424F33468B096FCF452AE0505A185905CC2414D44437118630839B88",
INIT_07 => X"588C732074A68D5AB4EB180717FF513FC52691924098712CE481FDC201D43C1A",
INIT_08 => X"0016053F180A1286A4ED1BC18840C320000055FE91AA545CBA4DE1D17992D9BE",
INIT_09 => X"2D1A4D8105B734723041008100486100601EDE1DE46431138DFD404CB4022595",
INIT_0A => X"A131112C0D15C901B2122309204C28B67061E81A8920C8D3CF8014007902DA6B",
INIT_0B => X"AD5C3402488888E5126BA350B27C092E63D18C9C500577EEA33EF24C09B42464",
INIT_0C => X"096B80D6B80B6B80F6B8096B80F6B80B6B80D15C04B5C07AD50C94020D233107",
INIT_0D => X"8948020D829FA454104132252011E542387F810480C840C383751EF5606E0178",
INIT_0E => X"000200CA7FE0627FD25845E42151648F854480A042512028100A8C38280AA04C",
INIT_0F => X"D06101C55DE5E3E3C017E37FC3E0017C3F8817E37FC3E0017C3F900040241001",
INIT_10 => X"6CD381C0118797FE0817EA7FC3E0017C3F8817EA7FC3E0017C3F9900DFFFDE15",
INIT_11 => X"F800DFFFBE34F00C0270F3F55F1F8007FDBEBE25E0700463E1FF2C7E014FF7BE",
INIT_12 => X"C5DEF64EC090626FE40140459759173BBD6EF37D523E6030061341F07FD571F8",
INIT_13 => X"0C4DFE2A6FE2AC3082637F281BFFFC07E00007E07F7253D38337D1D6184131BF",
INIT_14 => X"4F4F8397FFA0F0E06101C53E76D3D3E884FDDDA8381C0098E5FD92BBDFC8D812",
INIT_15 => X"19074FA36FDF58DBF81C072540049707E0FEF313D3E03BFFF61478040570EFD5",
INIT_16 => X"8CA02ACA00C50850182309444D248204201040FC190054A2110B8ACC483204A1",
INIT_17 => X"0A128CA0284A2280A1288A128CA2284A0288A1288A3284A228CA0288A1280A32",
INIT_18 => X"A228CA0284A3280A3288A1288A3280A2284A028CA2284A2284A028CA0280A328",
INIT_19 => X"F6A1850E1892596D34924B2DA6A84A2284A1288A1280A3280A1288A0284A2284",
INIT_1A => X"7DF7DF7DF7CBFBFE7EFEEE79E79EFAF3F51EB769CFEF73B6FFE74FC2400DB6DB",
INIT_1B => X"EEF77BBDDEEF77BBDDEEF77DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF",
INIT_1C => X"FFC27F6BDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDD",
INIT_1D => X"55D2E955FFF7FFC0000000000000000000000000000000000000000000000200",
INIT_1E => X"EFAA84001FF5D043FEAA5D04020AA002AAAABA555140155087FFFFEF00042AB5",
INIT_1F => X"1550800001FF5D00001555D2E975FF5D5568B555D7BD5545FFD540155FF843FF",
INIT_20 => X"FF45A2FFC0000AAAE974AAFFFFEAA10F7D57FEAA557BE8B45A2D5555EFAAD540",
INIT_21 => X"401555D04174AA002A80010FFAE975FFAA80001EF002AAAABAF7D168A10A2D17",
INIT_22 => X"EBFEBA555542000A28028BFFF7803DF55FFAEBFE005D2EAAB45557BD55555555",
INIT_23 => X"517DF55082E974BA087FE8B55552E955EF5D7FEAA105555421EFFFD568AAA002",
INIT_24 => X"00000000000000145FF842AAAAA2AA800BA5D51555EF002AA8BFFAAAA820AA5D",
INIT_25 => X"007FFFFFF1C042FB7D492A955C7F7FBC00000000000000000000000000000000",
INIT_26 => X"5E3DB45145E3803AFEFA284051D755003DE92410F42092142E28ABA5D5B4516D",
INIT_27 => X"6DBEDF575FFAADF42155082E851C75D0E02145492E955C75D5F6DB55497BD554",
INIT_28 => X"ABAF7D16DA28A2DB7AF7DB6FBC7028A2AA95492FFFFE8A38EBD57DE824975EAB",
INIT_29 => X"FB45557BD5555415F45145490A124BA002080010FFA4955C7BE8E021C71C0A2D",
INIT_2A => X"451D7EBD16FAAA002ABFEAA555F42000E2AAA8BEFE3843AF55E3AABFE105520A",
INIT_2B => X"4821D7F68E07082495B7FF7D082E954AA087FEDB7D5D2A155D7157BEFA38555F",
INIT_2C => X"0000000000000000000000000000002145F7802AABAA2A480092415B505D7142",
INIT_2D => X"52CAAAAA5D7FD75EF087BFDFEF5D003DFEF002E95555F7FDC000000000000000",
INIT_2E => X"5D7BFDF45007FD7555A2F9D5555A2802ABFFAA841754555043FE10082A820005",
INIT_2F => X"AAAD57DE1000516ABFFFFFBD75FFAAFFC0145002895545552E80145002E95545",
INIT_30 => X"45F7AE821455D2CBFEAAFFD17FEAAAAFFEABFFF7FFD54BAA2AA95410F7FDEAAB",
INIT_31 => X"B45AAAABFE0009043FF555D7BD55550879D5555002E820BA080400010FF80175",
INIT_32 => X"75455D7DFFEBA5D7BD5545A2D57DEAA002EBDEAA557BC0000AAA8A8BEFA28028",
INIT_33 => X"02010007FC0155550222955FFAC97400087FFFFFF002E954AA087BFFFFF5D2E9",
INIT_34 => X"000000000000000000000000000000000000000000000000155F7802AAAAAA80",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000003000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B0061A258A2840112C03002C180004003220200403302301C0381A0086",
INIT_01 => X"860041C83839484C00A100000052024841000000090800090210010000510204",
INIT_02 => X"080108200C1000004464080400C0080100000000010432400800800009882050",
INIT_03 => X"040001008C2340D0800208624200002183800584488000103080010C08C10000",
INIT_04 => X"00101610A029B08400044800000000040008102A040810040400900500001800",
INIT_05 => X"02800000400C830934E4A0002900404400820000000A00824004084011200A00",
INIT_06 => X"14C8874C884D0C024608680210C11F8010122100880802800308010000829400",
INIT_07 => X"060800002430200004611000508184803A0900224000200008818028C04883E1",
INIT_08 => X"4041FE80E009024260240010608000000000043E040000488000201400008810",
INIT_09 => X"0002447E041B112020208010404029006FE0B081003204502000002068621191",
INIT_0A => X"35E5148B0D916BBE39049191200000200441048108000220002FC5FA60000148",
INIT_0B => X"5358BF12E88D1000022808801A112D1443142A815440600083FE9AA300100281",
INIT_0C => X"C1416C1416C5416C5416C3416C3416C7416C500B60A0B60AD40E34104C093904",
INIT_0D => X"8C03403C440C054048850A300A8480009A0020865AE4ECB11B441A105B05B016",
INIT_0E => X"00000031001E4800022100321489214001A742D3A368D1B4686D100234B44242",
INIT_0F => X"00000000000AB800302008000000014000602008000000014000674000260000",
INIT_10 => X"0000000000000241E020010000000140006020010000000140006A8400000000",
INIT_11 => X"028400000000000000000003C00052000200000000000000000CD00184000800",
INIT_12 => X"30000800000000049A48184000A0400000010000000000000000000048028C00",
INIT_13 => X"0000918480010000000024C9E000000000000000000FF0006440200000000012",
INIT_14 => X"C000602800400000000000000BB000112B0020000000000000007E0000010000",
INIT_15 => X"02A0005000202500010000000000000000104CF000198000000000000000000F",
INIT_16 => X"4AD2B46D180684E8402440044C24A30819020603E0A20640C8400010218432A0",
INIT_17 => X"2D1B4ED3B4AD0B42D1B4ED2B42D0B46D1B4ED2B42D1B46D3B4AD2B42D1B46D2B",
INIT_18 => X"D1B42D0B46D2B4AD1B46D0B4AD3B4ED0B46D1B4AD2B4ED1B42D0B4ED3B4ED0B4",
INIT_19 => X"F8840000331C618E38E38C31C7346D3B4AD3B46D0B42D3B4ED2B42D1B42D2B4E",
INIT_1A => X"1C71C71C71CEDBB676F66EFBEFBEFAF99CFEF179CFF1FE1E9F52AFF9BFAFBE7B",
INIT_1B => X"FE7F3F9FCFE7F3F9FCFE7F1C71C71C71C71C71C71C71C71C71C71C71C71C71C7",
INIT_1C => X"FFE43591FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"05D2EBDF55557FC0000000000000000000000000000000000000000000030200",
INIT_1E => X"55087FFFFEF00042AB555D2E955FFF7FFC21EFF7D17DEAA5D2AAAAAA5D557DE1",
INIT_1F => X"0AA002A82145555542010FF803DEAA5D5568BEF5D042AA10A2AAAAABA5551401",
INIT_20 => X"20BA00557DF455D7BFFEAA555540155FF843FFEFAA84001FF5D043FEAA5D0002",
INIT_21 => X"001FF5D00001555D2E975FF5D5568B555D7BD5545FFD568AAA5D00154AAAAD14",
INIT_22 => X"5555EFAAD540155080000000F7843FF55007FFDEAAA284020BAAAD168BFF0800",
INIT_23 => X"51401EFF7842AA00FF8417545AAAEBFE10FFFFEAA10F7D57FEAA557BE8B45A2D",
INIT_24 => X"0000000000002AABAF7D168A10A2D17FF45A2FFC0000AAAE974AAFFFFC21EF55",
INIT_25 => X"5520ADA92495B7AE10412EBFF45497FC00000000000000000000000000000000",
INIT_26 => X"0AAAAA8ABA5D5B4516D007FFFFFF1C042FB7D492A955C7F7FBC71EFFFD57FE82",
INIT_27 => X"D755003DE92410E02092140E0716D415F47000F78A3DE92415F6ABD7490A28A1",
INIT_28 => X"A92550A104AABED1470AA005F78F7D497FFFE925D5B45145E3803AFEFA284051",
INIT_29 => X"20BAA2DB68BC7140E051C75D0E02145492E955C75D5F6DB55497BD5545E3DB6A",
INIT_2A => X"7DE824975EAB6DBEDF575FFAADF42155082E87038FF8038F6D1C7BF8EAAAA800",
INIT_2B => X"A95492FFFFC71EF415F471C7FF8428A00E38412545AAAE3FE10A3FBE8A38EBD5",
INIT_2C => X"000000000000000000000000000002DABAF7D16DA28A2DB7AF7DB6FBC7028A2A",
INIT_2D => X"7FDD55EFF7D57DE005D003DE00007FEAA10002ABFF450079C000000000000000",
INIT_2E => X"087BE8B45082EAAA10A2A8AAAAA5D7FD75EF087BFDFEF5D003DFEF002E95555F",
INIT_2F => X"5A2802ABFFAA841754555043FE10082A82000552C955FF007BD5410FFAABFE00",
INIT_30 => X"45007FD7555A2F9EAA005D2A820AAF7D5574AA087BEABEF007FFDE00557DD555",
INIT_31 => X"BFF557BE8ABAA284020BAA2FBEAB55552C95545552E80145002E955455D7BFDF",
INIT_32 => X"FE10A2F9EAABAAAD57DE1000516ABFFFFFBD75FFAAFFC01450028974BAFF842A",
INIT_33 => X"EABFFF7FFD54BAA2AA95410F7FDD55EF007BD5555F7802AA10AA8000145AAAEB",
INIT_34 => X"00000000000000000000000000000000000000000000003FEAAFFD17FEAAAAFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000002400000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0048201002842002C02450018800002300500030B313300C418992002",
INIT_01 => X"A34009C23838684D1C20E0000E11426840000000080000080200080000110200",
INIT_02 => X"4801082048100000446558040080000041000000000622400800000009000010",
INIT_03 => X"040001818CA144D0842248424210812103000480088000003080014688800000",
INIT_04 => X"000012002041900000048000000000040088322944200C850001940400301800",
INIT_05 => X"0200000040084000284000204104004402000025000800065004207030320800",
INIT_06 => X"108017080149000246086A2A1468004012120004440812D40120008200829001",
INIT_07 => X"2408000024302040846810005281848003494020400031240C8C8218E06A0009",
INIT_08 => X"4040050001090242602C0418408000000000243E0408104C8000201540008810",
INIT_09 => X"00024401041B132820000001424069004000B204636009104A0101226A422104",
INIT_0A => X"80049800A0281400300B0210200008B206639389480046240068180262000048",
INIT_0B => X"41401C1081811C44D22A18841616004118004482040448011800004D49340082",
INIT_0C => X"00192001920019200192041920419204192060C9010C90100008040008012101",
INIT_0D => X"48A000880144434A001001228000803198003604004048294008C40C483480D2",
INIT_0E => X"0000002160006000100000200811020805000480004000220108000060000800",
INIT_0F => X"09864038A2881210382000000001E003E0582000000001E003E0422834240000",
INIT_10 => X"0000160700706901982000000001E003E0582000000001E003E04E8400000000",
INIT_11 => X"0684000000000330C00F0C8210807200000000000581C01C1C809201C4000000",
INIT_12 => X"29D000000C2419121028C00020A2400000000000080082C180603A0E003A0904",
INIT_13 => X"8322414E800000432118908DF8000000061E001FC00C10207740000021908C48",
INIT_14 => X"40806BB800000009864038C14810201BAB000000026130071A80613A00000184",
INIT_15 => X"840080546520350000600812058100F81C018890201BBA0000008239020F1108",
INIT_16 => X"04812208033400C0022140404D268624B210040004A08400000044222900320C",
INIT_17 => X"0832048120481204822008020080204832048120480200802008020081204812",
INIT_18 => X"802008020C812048020080200812048120080200802048120483200802008020",
INIT_19 => X"0221054A2C208200010410400020880200812048120C80200802008120C81200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFD3B3D800000000000000000000000000000000000000000000000000000000",
INIT_1D => X"5AA8017410555540000000000000000000000000000000000000000000000200",
INIT_1E => X"AA5D2AAAAAA5D557DE105D2EBDF55557FFDE00557BEAABAA2AEAABEFF7801555",
INIT_1F => X"5FFF7FFD5555557BEABFFF7FBEAAAAAAD157555AA803FEBA5555421EFF7D17DE",
INIT_20 => X"DFEFAA80000BAAAAA820BAA2802AABA555140155087FFFFEF00042AB555D2E95",
INIT_21 => X"02145555542010FF803DEAA5D5568BEF5D042AA10A2AA955EFF7FFD5400F7FFF",
INIT_22 => X"43FEAA5D00020AA002ABDEBA5D7FE8A000004154BAF780001EFAAAAA8B450000",
INIT_23 => X"2AAABFF5551421FFAAD157545AAD5555EF557FC0155FF843FFEFAA84001FF5D0",
INIT_24 => X"00000000000028AAA5D00154AAAAD1420BA00557DF455D7BFFEAA5555575455D",
INIT_25 => X"AAA0A8BC7EB8417555AA84104385D55400000000000000000000000000000000",
INIT_26 => X"A4155471EFFFD57FE825520ADA92495B7AE10412EBFF45497FFFE385D71E8AAA",
INIT_27 => X"FF1C042FB7D492A955C7F7FBD056D5D75EABC7FFF5EAAAABEDF5257DAA8438EB",
INIT_28 => X"5EFEBFFD2400EBFBFAFEFAA80070BAA2A0870BAAA8028ABA5D5B4516D007FFFF",
INIT_29 => X"01D7AAA0AFB6D1C040716D415F47000F78A3DE92415F6ABD7490A28A10AAAA92",
INIT_2A => X"3AFEFA284051D755003DE92410E02092140E3DE924171E8A281C0E10482F7840",
INIT_2B => X"FFFE925D5B525454124AFBC74955421EFA2DF5557DAAD5D05EF0175C5145E380",
INIT_2C => X"000000000000000000000000000002AA92550A104AABED1470AA005F78F7D497",
INIT_2D => X"079FFEAA5D5568ABAA2842AB55A28015545A284000BA5D534000000000000000",
INIT_2E => X"F7FBC01EFA2842AABA0857555EFF7D57DE005D003DE00007FEAA10002ABFF450",
INIT_2F => X"A5D7FD75EF087BFDFEF5D003DFEF002E95555F7FDC01EF55556AB55F7D56AABA",
INIT_30 => X"45082EAAA10A2A8801FFA2FFC2000A2FFEABFFAA84174BAAA80174AAAA862AAA",
INIT_31 => X"AAA552A80010F78000145AA843DFEF5D02155FF007BD5410FFAABFE00087BE8B",
INIT_32 => X"21FF085755555A2802ABFFAA841754555043FE10082A82000552CBFE10085168",
INIT_33 => X"574AA087BEABEF007FFDE00557DC014500003FF450051401FFA2FBD55EFAAD54",
INIT_34 => X"00000000000000000000000000000000000000000000002AA005D2A820AAF7D5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"A14008420008204D042100000212026840000000180800080200090048510204",
INIT_02 => X"080108000090000004655C040080000051000000000402400800000009000010",
INIT_03 => X"00000100803008D0842240024210810003800584488000103080894288800000",
INIT_04 => X"00009610A028B084000440C0040000040088323244280C950400808500321800",
INIT_05 => X"42800080400C8A09306420202804400402800035200A00020204287001114A00",
INIT_06 => X"14C8864C8849880002486800142BFF001292214444081254002801A200821400",
INIT_07 => X"004800002430204084281000D281040001182020400031241C0D80000041BFE9",
INIT_08 => X"444005000108020220240010048000000000043E0408104C8000000100008810",
INIT_09 => X"0812040105191100200081130210ED104008A285617205D02A01010141225091",
INIT_0A => X"8004C8252291490039039390200008B20E230008280040088040100240008061",
INIT_0B => X"40013C128BC95C44522A00241204094008442681100448000800826F49240001",
INIT_0C => X"0408000080000800008000080000800008000440020400229548040008012125",
INIT_0D => X"401140BC4028430108150900408590109A00209642E46CA00240460400200440",
INIT_0E => X"080410010000200002210A320C89000005A142D0A16850B6294D100234201242",
INIT_0F => X"2F9EC00000800008100020003C1FE00020080020003C1FE00020044014260082",
INIT_10 => X"132C7E3F00000100080020003C1FE00020080020003C1FE000200880000081EA",
INIT_11 => X"0080000081CB0FF3C000008000201000010001DA1F8FC0000080110080000010",
INIT_12 => X"040000B0BE6C00020040580040200000001004832CC19FCF81E0000000100002",
INIT_13 => X"80004020000C31CF60001000000007F01FFE00004000300420000618E7B00008",
INIT_14 => X"C0102000000F151F9EC0000040300401000200D547E3F00000800080001617AD",
INIT_15 => X"02A020100000822406E1B95A3F83000000008030040100000BAB87FB00000100",
INIT_16 => X"46D1B66D1A368C68D26000544D26A504AB120400222206404840001101843000",
INIT_17 => X"2D1B46D1B46D1B46D1B46D1B46D1B42D0B42D0B42D0B42D0B42D0B42D1B46D1B",
INIT_18 => X"D1B46D1B42D0B42D0B42D0B42D1B46D1B46D1B46D1B42D0B42D0B42D0B42D0B4",
INIT_19 => X"20840442200000000000000000346D1B46D0B42D0B42D0B42D0B42D1B46D1B46",
INIT_1A => X"3CF3CF3CF3DBF91E66C6FAD96D965201F4C251414A87D78AF421448BE28F3AEB",
INIT_1B => X"3E1F0F87C3E1F0F87C3E1F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"FFD160B27C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C",
INIT_1D => X"AFFFFC2000557FC0000000000000000000000000000000000000000000000200",
INIT_1E => X"BAA2AEAABEFF78015555AA80174105555420000000021EFAA843DE00F7803FEB",
INIT_1F => X"F55557FD54AAA2AA955FF00043DE005504175FF08514014555557DE00557BEAA",
INIT_20 => X"DF45FFD17DFFFFFD56AA00557FC21EFF7D17DEAA5D2AAAAAA5D557DE105D2EBD",
INIT_21 => X"55555557BEABFFF7FBEAAAAAAD157555AA803FEBA55556ABFFA280154BAFF803",
INIT_22 => X"42AB555D2E955FFF7FFD5410002AAAAAAA2D57DF450004154BA087BEAAAAF7D5",
INIT_23 => X"843DE1008556AA00A28028B55FFD1555EFA2802AABA555140155087FFFFEF000",
INIT_24 => X"000000000000155EFF7FFD5400F7FFFDFEFAA80000BAAAAA820BAA280000AAA2",
INIT_25 => X"A2803AE38FF843DEBAEBFFC20285D75C00000000000000000000000000000000",
INIT_26 => X"55D5F7FE385D71E8AAAAAA0A8BC7EB8417555AA84104385D5542038000A001C7",
INIT_27 => X"92495B7AE10412EBFF45497FD24BAA2AA955C708003FE285D00155FF00554515",
INIT_28 => X"BEFA28E124AAF7843AF7DEBDB78FFFE3DF6DA284175C71EFFFD57FE825520ADA",
INIT_29 => X"04920875EAA82F7DB5056D5D75EABC7FFF5EAAAABEDF5257DAA8438EBA415568",
INIT_2A => X"4516D007FFFFFF1C042FB7D492A955C7F7FBD54380020ADA82BED57DF4508041",
INIT_2B => X"0870BAAA80070BAA2803DE00005F68A10BE802DB55E3DB555FFF68028ABA5D5B",
INIT_2C => X"00000000000000000000000000000125EFEBFFD2400EBFBFAFEFAA80070BAA2A",
INIT_2D => X"D53420BA082E82155AA802AAAAFF803DEBAAAFBC20BA55514000000000000000",
INIT_2E => X"5D04175EF0855575455D7BFFEAA5D5568ABAA2842AB55A28015545A284000BA5",
INIT_2F => X"FF7D57DE005D003DE00007FEAA10002ABFF450079C20BAAAAE9754500043DEBA",
INIT_30 => X"EFA2842AABA085768BFFA2AE820AAFF802ABEFAAFFEABEFAAFFFDEAA0051555E",
INIT_31 => X"E10F7D17FF5500000001008516AA10FFFFC01EF55556AB55F7D56AABAF7FBC01",
INIT_32 => X"75EFF7842AAAA5D7FD75EF087BFDFEF5D003DFEF002E95555F7FDD74BA08043D",
INIT_33 => X"EABFFAA84174BAAA80174AAAA86174AAAA843DE00087FE8A00F7843FF45AAFFD",
INIT_34 => X"0000000000000000000000000000000000000000000000001FFA2FFC2000A2FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000001000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"A1400802000020490000000000000240413C0A61590001D90213C90008510204",
INIT_02 => X"680108200010000054655C040080000041000000010402400800800009082011",
INIT_03 => X"00040100800020D0842240124210810043800504488000103081894288800000",
INIT_04 => X"00001410A00AA084000400C0060000040088323044201C850020820400101880",
INIT_05 => X"0200020040048A09202420000C00410402000025000800020804207000100800",
INIT_06 => X"10488704884D080202086A0A3429004012120004DC08125400A0008300821000",
INIT_07 => X"000800002C30204084381000128104000100002040003164040D800000400009",
INIT_08 => X"0440050003080202202400100080000000000C3E0408104C8000102300008810",
INIT_09 => X"4810240104111104200080120210A5104000A204615201500801010000AA10C0",
INIT_0A => X"81F525A82804010009029290200008B202238008080240000040100242048025",
INIT_0B => X"00A1141002C91844522A0004120488000800028000044000080020AF09240010",
INIT_0C => X"0408104081000810408100081040810008104040800408208040000008010121",
INIT_0D => X"4201E0B4000803200C150108008490809A002192462424202200440404204041",
INIT_0E => X"0804100160006000120002120499020A04A14650A32851962965190014200240",
INIT_0F => X"000000000080A200100021000000014020080021000000014020000014260082",
INIT_10 => X"0000000000000340080028000000014020080028000000014020008000008000",
INIT_11 => X"008000008000000000000081500010000100800000000000008C100080000012",
INIT_12 => X"05D0000880000006800058000020000000000005000000000000000048100100",
INIT_13 => X"0000D02E8040200000003401F80004000000000040026000274000900000001A",
INIT_14 => X"800023B8000030000000000042A00009AB00008800000000008012BA01001000",
INIT_15 => X"00A000106520350000040100000000000010C0200009BA000200000000000105",
INIT_16 => X"465196651B328CA8D26540544924272EB91004002022024048400000098030A0",
INIT_17 => X"6509425094250942509425094250942509425094250942509425094251946519",
INIT_18 => X"5094250942509425094250942519465194651946519465194651946519465194",
INIT_19 => X"2A05404808000000000000000014651946519465194651946519465094250942",
INIT_1A => X"69A69A69A68945B080201C92410480ABD102E689999E91BCD151200C30AE1C71",
INIT_1B => X"341A0D068341A0D068341A28A28A28A28A28A28A28A28A28A28A28A28A28A69A",
INIT_1C => X"FFC5B52068349A4D068341A0D269341A0D269341A0D068349A4D068349A4D068",
INIT_1D => X"0F7D17FFFFAAAE800000000000000000000000000000000000000000000003FF",
INIT_1E => X"EFAA843DE00F7803FEBAFFFFC2000557FEABEFA2D1400AA5D2AAAA00F7FFEAA1",
INIT_1F => X"4105555421EFF78028BEF5D003DFEFF7FFE8ABAF7802ABEFAAAE820000000021",
INIT_20 => X"AB45557BC0155007FFDEBAAA843DE00557BEAABAA2AEAABEFF78015555AA8017",
INIT_21 => X"154AAA2AA955FF00043DE005504175FF0851401455555555EFA2FBC01FFF7AAA",
INIT_22 => X"57DE105D2EBDF55557FFDE00552A974AAA2843DEAA5D2A820BA000428AAAAA84",
INIT_23 => X"517FFEFAAAEBDF45FFAEA8ABAF7D1400BAAAAE821EFF7D17DEAA5D2AAAAAA5D5",
INIT_24 => X"0000000000002ABFFA280154BAFF803DF45FFD17DFFFFFD56AA00557FC201000",
INIT_25 => X"4120ADA38E3F1EFA28F7DF7DFD7A2A4800000000000000000000000000000000",
INIT_26 => X"7A2A482038000A001C7A2803AE38FF843DEBAEBFFC20285D75EFBC7A2DB40082",
INIT_27 => X"C7EB8417555AA84104385D55421C7FF8028BEF41003FFD7F7F1EDA82F78E2DBD",
INIT_28 => X"5C7A2FBC51EFEBA0A8B6D5571C716D1475FFEAAA28E3FE385D71E8AAAAAA0A8B",
INIT_29 => X"50AA1C0428ABAB68E124BAA2AA955C708003FE285D00155FF0055451555D5F57",
INIT_2A => X"7FE825520ADA92495B7AE10412EBFF45497FFFE105D2E97482AA8038EAA412E8",
INIT_2B => X"F6DA284175C001000557FFEFB6A0BFF55F7AEAAA82FFDF40092B6A4871EFFFD5",
INIT_2C => X"0000000000000000000000000000028BEFA28E124AAF7843AF7DEBDB78FFFE3D",
INIT_2D => X"5517DF55A2FBC201008003DEAAA2D57FEAAF7FBFDF45AA800000000000000000",
INIT_2E => X"FFD57FE00FFAABFF45AA80020BA082E82155AA802AAAAFF803DEBAAAFBC20BA5",
INIT_2F => X"A5D5568ABAA2842AB55A28015545A284000BA5D5340145F78028BFF08003DF45",
INIT_30 => X"EF0855575455D7BD5555A2FBD75FFA2842ABFF5555575FF55557FEAAA2AABFEA",
INIT_31 => X"400A2802AABA002A954AA5D0028ABAF7AA820BAAAAE9754500043DEBA5D04175",
INIT_32 => X"2010FF80155EFF7D57DE005D003DE00007FEAA10002ABFF450079FFE005D2A97",
INIT_33 => X"2ABEFAAFFEABEFAAFFFDEAA00514200008517DFEFFF803FF45FFAAA8A00F7FBC",
INIT_34 => X"000000000000000000000000000000000000000000000028BFFA2AE820AAFF80",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000002000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033022000000180006",
INIT_01 => X"0000098218302849180060000C00424040000000080000080200090008510200",
INIT_02 => X"0801080200100000044008000080000041000000002002400800000009008010",
INIT_03 => X"0001000004000040000202000000000803006400088000003080040008C10000",
INIT_04 => X"0000100022008000000C08C00C00000400201830040000040000000400001820",
INIT_05 => X"0200000040000000248080210044000400000000000800000004000010000800",
INIT_06 => X"100007000049000202086A080000004010100000880800001000000030829000",
INIT_07 => X"000800002420000004201000128100000300002040003124040D802040400009",
INIT_08 => X"040005000108020220240020008000000000043E000000488000000100008811",
INIT_09 => X"0810040105111000202000024010A51040088080000000110000002000020084",
INIT_0A => X"040000000000010000040010200008B202230480080002000000100240008021",
INIT_0B => X"40003C020AC04400022808001000014000040088140000000000828000000820",
INIT_0C => X"0040004400044000040000400044000440000400002000221048840009012124",
INIT_0D => X"0002A00800000100440000000800800018002000008000800040022000000400",
INIT_0E => X"0804100100002000100002001001024800020001000080004000000800904000",
INIT_0F => X"000000000000A000102008000000014000082008000000014000000000240082",
INIT_10 => X"0000000000000240082001000000014000082001000000014000028000000000",
INIT_11 => X"028000000000000000000001400012000200000000000000000C100084000800",
INIT_12 => X"0000080000000004800000400020400000010000000000000000000048000000",
INIT_13 => X"0000900000010000000024080000000000000000000250002000200000000012",
INIT_14 => X"4000200000400000000000000290000100002000000000000000120000010000",
INIT_15 => X"0000001000000000010000000000000000104010000100000000000000000005",
INIT_16 => X"0000000001400080002100544924002A000004000020000080000000010032A0",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100400000000",
INIT_18 => X"0000000000000000000000000010040100401004010040100401004010040100",
INIT_19 => X"02A1410808000000000000000000000000000000000000000000000000000000",
INIT_1A => X"145145145146AB2A0CCC2A28A28A7AA0CDF0D1215281FC1A72E24C28E921AAA9",
INIT_1B => X"CA6532994CA6532994CA65145145145145145145145145145145145145145145",
INIT_1C => X"FFD9C63B95CA6532994CA6532B95CAE572994CA6532994CAE572B95CA6532994",
INIT_1D => X"FAAD1555FFF78400000000000000000000000000000000000000000000000200",
INIT_1E => X"AA5D2AAAA00F7FFEAA10F7D17FFFFAAAE801FF08557DF4555516AA00007BEABE",
INIT_1F => X"000557FC0010AAD57FF45A2D56AA0000043FFEFA2FFFDE1008556ABEFA2D1400",
INIT_20 => X"DEAA007FEAB45AAAE800AAF784020000000021EFAA843DE00F7803FEBAFFFFC2",
INIT_21 => X"421EFF78028BEF5D003DFEFF7FFE8ABAF7802ABEFAAAEA8BFF5D0415400F7FBF",
INIT_22 => X"015555AA80174105555401FF5D0415555557BFDFEF00517DE00A28028B450855",
INIT_23 => X"FFD7555AAD56AB45A2AE800AA5D7FFDEBAF7AEBDE00557BEAABAA2AEAABEFF78",
INIT_24 => X"000000000000155EFA2FBC01FFF7AAAAB45557BC0155007FFDEBAAA8417410AA",
INIT_25 => X"55556AA381C75EABEFBED1575C7E380000000000000000000000000000000000",
INIT_26 => X"81C516FBC7A2DB400824120ADA38E3F1EFA28F7DF7DFD7A2A4801EF085F7AF6D",
INIT_27 => X"38FF843DEBAEBFFC20285D75C0010AADF7AF6DB6D56FA3814003AFFFA2F1F8E3",
INIT_28 => X"BEF550412428F7F5FDE920875E8B45BEA0850BAE38002038000A001C7A2803AE",
INIT_29 => X"8E10AA802FB450851421C7FF8028BEF41003FFD7F7F1EDA82F78E2DBD7A2A4AD",
INIT_2A => X"E8AAAAAA0A8BC7EB8417555AA84104385D55401C75504125455575FAFD714557",
INIT_2B => X"5FFEAAA28E10438AAF5D2545BED56FB45BEA082082557BF8EBAF7AABFE385D71",
INIT_2C => X"00000000000000000000000000000175C7A2FBC51EFEBA0A8B6D5571C716D147",
INIT_2D => X"A80021FF007BE8BFF5D516AABA5D5568BEFF7D157555AA800000000000000000",
INIT_2E => X"5D002ABFFA2D16AAAA55517DF55A2FBC201008003DEAAA2D57FEAAF7FBFDF45A",
INIT_2F => X"A082E82155AA802AAAAFF803DEBAAAFBC20BA555140010AAFFE8BFFFFD17DEBA",
INIT_30 => X"00FFAABFF45AA803FFEF5500020BAFFD17DE10005568B55FF80154BAA280020B",
INIT_31 => X"1555D556AB555D5568A00AA843FF55085140145F78028BFF08003DF45FFD57FE",
INIT_32 => X"AAAAF7AABFEAA5D5568ABAA2842AB55A28015545A284000BA5D5342145550402",
INIT_33 => X"2ABFF5555575FF55557FEAAA2AA800AAAAD142155F7D57DF45FF8002010557FE",
INIT_34 => X"000000000000000000000000000000000000000000000015555A2FBD75FFA284",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000023FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B830084C1820E0000C36424840000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"000406A492E6E440842254D002108153422004800880000030C0315688C00006",
INIT_04 => X"00001201200090001205400000000094108C322644240C840008030440111800",
INIT_05 => X"222000444008010028404002A002009402400025080880000C04223000170900",
INIT_06 => X"12801628014B0B000A086CA6556800C012121004540816544522008200821100",
INIT_07 => X"1C08320054B624408428100094ADD080011721A04000316C140CA1A8A1F90019",
INIT_08 => X"00140500090B02C2E0EC04D1C08000000000647E858A104C920C81A5011088A6",
INIT_09 => X"40002481041F165820000101024061004004800567603592A801014C46426011",
INIT_0A => X"8404002020000101B0070310200008B60A23A51B28024CE24E40100260040004",
INIT_0B => X"2800340208811865D22BB384100E01090805A495100400050800E24D49A424C5",
INIT_0C => X"0C72A0872A0C72A0872A0C72A0C72A0872A0C595043950421400800009010104",
INIT_0D => X"4290A088812203360410110A400085539800210404C048CAC040464D28014405",
INIT_0E => X"0804101160006000101004A01811064B050204810240812241280D00200A0804",
INIT_0F => X"6D0141B0482A01AAEC3602330CD2A02952DC3502330CB4A0318B414000240082",
INIT_10 => X"5B4551630144C0155C3502330CD2A02952DC3602330CB4A0318B5600C587149B",
INIT_11 => X"FE04E587083B6A51005956308D1E8202C436375908AA840AD4513437640F1524",
INIT_12 => X"E020C67062F47B2872400044959BC42B1060F0D036B80B548523136C158878D8",
INIT_13 => X"8F0B27010A2699AAA3794392000D81852B0A050C224180062085134CD1719564",
INIT_14 => X"0AD57400C50500D94C8121713C02B555101C90705D71009604140C0418CE0C37",
INIT_15 => X"DC06A27C828E024D8C50965A40821568A06113801505010334AA73AA0666DAC2",
INIT_16 => X"04812048123408C0822040004C248604B2100400100084008001D0113920060C",
INIT_17 => X"4812048120481204812048120481204812048120481204812048120481204812",
INIT_18 => X"8020080200802008020080200812048120481204812048120481204812048120",
INIT_19 => X"00A0014200000000000000000020080200802008020080200802008020080200",
INIT_1A => X"4104104104140D220A4A380000002A80E900C4C1100830181621409C80210821",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000410",
INIT_1C => X"FFC1F83800000000000008040000000000000000000201000000000000000000",
INIT_1D => X"0F7842AA00002A80000000000000000000000000000000000000000000000200",
INIT_1E => X"4555516AA00007BEABEFAAD1555FFF784020AAF7D542155F7D1400AAF7FFFDE0",
INIT_1F => X"FFFAAAEA8ABAFFD17FEBAFFAA800AA007FFDFFFA28428A000000001FF08557DF",
INIT_20 => X"00AAF78028AAAFF84020AAFFFBEABEFA2D1400AA5D2AAAA00F7FFEAA10F7D17F",
INIT_21 => X"40010AAD57FF45A2D56AA0000043FFEFA2FFFDE1008556AB45555568A10A2FFC",
INIT_22 => X"03FEBAFFFFC2000557FC0155FFD1555FF0804000AA000428A10AAAA801EFFFD1",
INIT_23 => X"8428A10087FD7400552EBDFEFA2FBFFF550000020000000021EFAA843DE00F78",
INIT_24 => X"00000000000028BFF5D0415400F7FBFDEAA007FEAB45AAAE800AAF78428B45A2",
INIT_25 => X"E3DF450AAF7F1FDE38FF8A2DA101C2A800000000000000000000000000000000",
INIT_26 => X"01C0E001EF085F7AF6D55556AA381C75EABEFBED1575C7E380000BAF7DB4016D",
INIT_27 => X"38E3F1EFA28F7DF7DFD7A2A4AFABAFFDF7AE82F7AA870AA0071F8FFFBE842DA1",
INIT_28 => X"B455D5B68A28A2FFC20AAEB842DAAAE38A02082E3FBEFBC7A2DB400824120ADA",
INIT_29 => X"8A28AAA4801FFE3DF40010AADF7AF6DB6D56FA3814003AFFFA2F1F8E381C516D",
INIT_2A => X"001C7A2803AE38FF843DEBAEBFFC20285D75C2145F7DF525EF140A050AA1C002",
INIT_2B => X"0850BAE3802DB6DAA8A28A00007FD74284120BFFFFBEF1F8F7D080A02038000A",
INIT_2C => X"000000000000000000000000000002DBEF550412428F7F5FDE920875E8B45BEA",
INIT_2D => X"A80020BAFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE10552E8000000000000000",
INIT_2E => X"085568BEFF7803FE10552E821FF007BE8BFF5D516AABA5D5568BEFF7D157555A",
INIT_2F => X"5A2FBC201008003DEAAA2D57FEAAF7FBFDF45AA803FEBAFFFBEAA00F7AE974BA",
INIT_30 => X"FFA2D16AAAA55517DF55557FEAAAAA2FFC00AAAA803FEAAA2AA82000A2FFFDF5",
INIT_31 => X"1EF552E974BA550028ABAA280001FFAAFFC0010AAFFE8BFFFFD17DEBA5D002AB",
INIT_32 => X"ABFF082E820BA082E82155AA802AAAAFF803DEBAAAFBC20BA555142155F7FFC0",
INIT_33 => X"7DE10005568B55FF80154BAA2803FFFFA2AAAAA00007FD74BA08003DFFFFFD16",
INIT_34 => X"00000000000000000000000000000000000000000000003FFEF5500020BAFFD1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000002000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C048000C048400380000007026040000000080000088200002802153231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"210D050012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"0080100022408000060DE0000066630C70241827041000040800820480001AA4",
INIT_05 => X"0240000C400000003C808003E0C8001401000000040900020904004000070800",
INIT_06 => X"1800068000491300CF0969A421C0004018184000100804005784000130821200",
INIT_07 => X"7E8C53200CA4850224301807D1CB45900147E03040083124FC0CD0C8A1FF0019",
INIT_08 => X"0046050013081206A4A503A9E8C0812000001C7E11A24058B84D40E33992D98F",
INIT_09 => X"010004810491175C20000080000821004010C01086003C13E000004EDF020400",
INIT_0A => X"000000000000010000180018200408B27E234913E9000CFA09A8180248001000",
INIT_0B => X"ACA0141000800021826933E03662802B3001E09F000000023000000000000867",
INIT_0C => X"0832F0C32F0832F0832F0C32F0832F0832F0C197861978400000000208010100",
INIT_0D => X"05FA0201E7F3F01F40401C17E800C7F3380020000000006AE01180493C5BC1AF",
INIT_0E => X"000200F500002200004005002001408400000000000000000000053A4096F807",
INIT_0F => X"246FC1B17B2C53F2FC16691DB587201EDDF4162B1DB527201EDDC46070241001",
INIT_10 => X"2A67DF2A01D5CC9794162B1DB587201EDDF416691DB527201EDDD884272592D6",
INIT_11 => X"288007258E995D5A825DBA569F9FF02547068618CD3CC45B7863AE7EC00D4B12",
INIT_12 => X"F6208C6CCA5C33717461C045B5B182019473D19D7CCD856106F31A683621BDFC",
INIT_13 => X"866E2FB10A652CC8E3538BBA01624E51AA6C0469AC5493F5688532966471A9C5",
INIT_14 => X"4F9B740041E1F5759001B4AA1853E6D5144AA9C914C8608D2724A4C4118D992B",
INIT_15 => X"DE07EAD9825682D4A36C0B0B4B85112B2C4A05D3E6D5051893335EB0072AA85A",
INIT_16 => X"00000000008000000821000048260020000004001DC0800000010E7F70171401",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0100401004010040100401004000000000000000000000000000000000000000",
INIT_19 => X"2A21010808000000000000000000401004010040100401004010040100401004",
INIT_1A => X"4924924924890380800016A28A28802B10B83728C1111026C152A23010848658",
INIT_1B => X"6432190C86432190C86432082082082082082082082082082082082082082492",
INIT_1C => X"FFDE003AC964B2592C964B2592C964B2592C964B2592C964B2592C964B2592C9",
INIT_1D => X"5FFAA80155F78400000000000000000000000000000000000000000000000200",
INIT_1E => X"55F7D1400AAF7FFFDE00F7842AA00002AAAA10FF8002155F7FFC200008041755",
INIT_1F => X"5FFF7842AB55080000145557FE8AAA080000155F7FFFDEAA0000020AAF7D5421",
INIT_20 => X"2000FF80020AAA2AAAABFF002E801FF08557DF4555516AA00007BEABEFAAD155",
INIT_21 => X"A8ABAFFD17FEBAFFAA800AA007FFDFFFA28428A00000028B4555043DFFFFFAE8",
INIT_22 => X"FEAA10F7D17FFFFAAAE80000A284174AAFF8428AAAFF8415545AAFBD7545F7AA",
INIT_23 => X"00000105D55400AA082A82155F7FFFDEAA08556ABEFA2D1400AA5D2AAAA00F7F",
INIT_24 => X"0000000000002AB45555568A10A2FFC00AAF78028AAAFF84020AAFFFBC215508",
INIT_25 => X"E3F5C000014041256DEBA487145F784000000000000000000000000000000000",
INIT_26 => X"2080E000BAF7DB4016DE3DF450AAF7F1FDE38FF8A2DA101C2AAFA00EB8E0516D",
INIT_27 => X"381C75EABEFBED1575C7E3802FB551C0E0516D417FEDA921C000017DEBF5FDE9",
INIT_28 => X"B55410A3FFC7F7A087000FF80070BAAAAAADBD70820801EF085F7AF6D55556AA",
INIT_29 => X"556DA2FBD7545F7AAAFABAFFDF7AE82F7AA870AA0071F8FFFBE842DA101C0E2D",
INIT_2A => X"400824120ADA38E3F1EFA28F7DF7DFD7A2A480000BE8A17482F78A28A92E3841",
INIT_2B => X"A02082E3FBC217D1C0E0500041554508208208017DF7F5FDE9208556FBC7A2DB",
INIT_2C => X"000000000000000000000000000002DB455D5B68A28A2FFC20AAEB842DAAAE38",
INIT_2D => X"52EBDE00AAAE975FFAAD1420005504001FFAA8015545F7800000000000000000",
INIT_2E => X"5504001FFAAD17DE00082E820BAFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE105",
INIT_2F => X"F007BE8BFF5D516AABA5D5568BEFF7D157555AA803DF45552E975EF007FFFE00",
INIT_30 => X"EFF7803FE10552EBDF45002EBFF55FF8017410FF84154BAAAAABFF450000021F",
INIT_31 => X"400F7AEA8A10A284175FFAAFBD5555F7AEBFEBAFFFBEAA00F7AE974BA085568B",
INIT_32 => X"DE1008517DF55A2FBC201008003DEAAA2D57FEAAF7FBFDF45AA8002000FFAE95",
INIT_33 => X"C00AAAA803FEAAA2AA82000A2FFC21EF552A954100851554000004021FFFFD17",
INIT_34 => X"00000000000000000000000000000000000000000000003DF55557FEAAAAA2FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00010100926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"0004122122029100100C00001200009C40A83A2044360C84190BAC04E0101820",
INIT_05 => X"027000004009050064C8C00104C10184034010250089C00EB004327064B60900",
INIT_06 => X"1B9416B94149000402086D42142800C012125804440812541027008230821380",
INIT_07 => X"0008320014B02848A4A8100015C55500057801A04000712C040CB1F880600009",
INIT_08 => X"005005000908020220E40170008042000000557E048A144C800590010000882D",
INIT_09 => X"0100250104B5310020000100020821004016CC1C616401910801010100CA2040",
INIT_0A => X"800000000000010192072310200028B6022346080802C0074AC0100259001004",
INIT_0B => X"A8201410008088C5D2288004120E802908800488000500050800404D49A42EB0",
INIT_0C => X"0400000000040000000000000040000000000000020000000000000008010102",
INIT_0D => X"4A02008000000360401021280800E400B800610C844848200028448400000000",
INIT_0E => X"000000086000600040D045E4195104D5854284A14250A12A512A880828984008",
INIT_0F => X"85D480949E07A80948354B6E68982167061037496E6838216706206810240000",
INIT_10 => X"652138E510B456587037496E689821670610354B6E6838216706220431961CA9",
INIT_11 => X"C2043196186A91674011CE61403562274AA49CD594CF00039C7C414B6509DA22",
INIT_12 => X"8A2E6A983014780CC8604040424A5323845932E620295879818170304B2F5002",
INIT_13 => X"8F019451654B9104A328665603148895D44E0251142B42A3D8B2A5C882519432",
INIT_14 => X"0AC5DC06A6C6A465AA0091482382B17614F2202858EE300991415B45CD530602",
INIT_15 => X"4000052E08DC8047F17D1C7C3C02128E587D6A02B17605A130A4E8BF00225885",
INIT_16 => X"84A1284A123508508220808048240604B2100C00022084809000D000393722A1",
INIT_17 => X"4A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A12",
INIT_18 => X"A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A128",
INIT_19 => X"F1228154000000000000000000284A1284A1284A1284A1284A1284A1284A1284",
INIT_1A => X"75D75D75D75FFAFEFEFEEEAAAAAAFBF3FC1FF77DDFE7EFBEFFE7CFC0044FBEFB",
INIT_1B => X"FAFD7EBF5FAFD7EBF5FAFD75D75D75D75D75D75D75D75D75D75D75D75D75D75D",
INIT_1C => X"FFC0003BF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5",
INIT_1D => X"F007FE8A00AAFBC0000000000000000000000000000000000000000000000200",
INIT_1E => X"55F7FFC2000080417555FFAA80155F7842AB55552E821FFFFD5555EF552ABDFE",
INIT_1F => X"A00002A821EF5D7BC21FFFFFBD55EFAAD1554BA00556AA00AAD16AA10FF80021",
INIT_20 => X"FF45A2AABFEBA082A975555D55420AAF7D542155F7D1400AAF7FFFDE00F7842A",
INIT_21 => X"EAB55080000145557FE8AAA080000155F7FFFDEAA00002AB45082A821EF5D557",
INIT_22 => X"BEABEFAAD1555FFF7842AABAA2FFE8BEF5D517FF455D554214500043DEBAAAFF",
INIT_23 => X"AABDF555D2E955EFA28428A10552EBFEAAAAD1401FF08557DF4555516AA00007",
INIT_24 => X"00000000000028B4555043DFFFFFAE82000FF80020AAA2AAAABFF002E80000AA",
INIT_25 => X"EBD5525C74124B8FC71C71EFA28AAF5C00000000000000000000000000000000",
INIT_26 => X"8AAD16FA00EB8E0516DE3F5C000014041256DEBA487145F78428B6D4120851FF",
INIT_27 => X"AAF7F1FDE38FF8A2DA101C2A871C74975C01FFEBF5D25EFA2D555482085F6FA2",
INIT_28 => X"B7D1C24851FF495F7FF55A2A0BFE921C2E9557D415B400BAF7DB4016DE3DF450",
INIT_29 => X"214508003FEAABEFFEFB551C0E0516D417FEDA921C000017DEBF5FDE92080E2A",
INIT_2A => X"7AF6D55556AA381C75EABEFBED1575C7E38028A82B6F1E8BFF495F78F7D49554",
INIT_2B => X"AADBD7082087000AAA4BFF7D5D20905C7AA842DA00492EBFEAABED1401EF085F",
INIT_2C => X"000000000000000000000000000002DB55410A3FFC7F7A087000FF80070BAAAA",
INIT_2D => X"78028BFF0004175EFA2D54214508042AB455D517DEBAA2D54000000000000000",
INIT_2E => X"AAD557410007BFDEAAA2D57DE00AAAE975FFAAD1420005504001FFAA8015545F",
INIT_2F => X"AFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE10552E975450051401EFA2D5421EF",
INIT_30 => X"FFAAD17DE00082EA8BFF5504175FF087BFFF45AA843FE005D2A955FF087BC20B",
INIT_31 => X"BFF087BEABEF00554215500003FEBAFFFBFDF45552E975EF007FFFE005504001",
INIT_32 => X"FEAAFFD5421FF007BE8BFF5D516AABA5D5568BEFF7D157555AA8028A00FFD16A",
INIT_33 => X"17410FF84154BAAAAABFF45000017410AA803DFEF550402155A2843FE00082AB",
INIT_34 => X"00000000000000000000000000000000000000000000003DF45002EBFF55FF80",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000033FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"000103A7A00904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000120122009000100C00000000000400A83A2044200C840000800400101820",
INIT_05 => X"020000004008010024C0C0010040000402000025000800020004207000100800",
INIT_06 => X"108016080149080002086807542800C012120004440812541020008230821000",
INIT_07 => X"4008120054B42850B42A100010ED1500010001A040003164040CF5E201400009",
INIT_08 => X"00400500090A020220A40A7000800000000014FE8508144C924080C100008801",
INIT_09 => X"0000040104111100200001000200210040008004616001910801010000422000",
INIT_0A => X"800000000000010190070310200008B202236D080802400002C0100240000000",
INIT_0B => X"0000141000800844522800041204000008000488000400000800004D49240820",
INIT_0C => X"0400004000000000000004000000000000004000000000000000000008010100",
INIT_0D => X"42020080000002204010010808008000B8002104044048200000440400000000",
INIT_0E => X"0000000000006000000000201811004005020481024081224128080820984000",
INIT_0F => X"CBA340480040A100A42008000161C140000420080001C1C14000032010240000",
INIT_10 => X"1A8A039600022260042001000161C140000420010001C1C140001604E8084341",
INIT_11 => X"1E04E8082580E2B8802201014800C220A21829A302F1C024010C001124020C8C",
INIT_12 => X"0024ACA60CA000048228404401004418012787124648157780120B8678C00080",
INIT_13 => X"00009001072D04730000241000CB1325E78E0186030240000083B60239800012",
INIT_14 => X"00001001EF6F4163C480481506800004000CFD55196CB012481812049495C194",
INIT_15 => X"40068248800108B8FB61A0401200845594965000000400568D0CFB7800550605",
INIT_16 => X"04812048123408408220000048240604B210040000008400800B0000090022A1",
INIT_17 => X"4812048120481204812048120481204812048120481204812048120481204812",
INIT_18 => X"8120481204812048120481204812048120481204812048120481204812048120",
INIT_19 => X"2820014000000000000000000020481204812048120481204812048120481204",
INIT_1A => X"3CF3CF3CF3CFFBBEEEEEFE79E79EFAABDDFAF369CB91FE1EF7D3AEBBDBAFBEFB",
INIT_1B => X"FE7F3F9FCFE7F3F9FCFE7F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"FFDFFFC1FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"AAAAEAAB45082E80000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFD5555EF552ABDFEF007FE8A00AAFBE8BEFA2D568ABA00003DF555555574A",
INIT_1F => X"155F78428AAA007FE8A1008002AABA555155400557BC2010557BEAB55552E821",
INIT_20 => X"FFFF082EBDEBAA2D1420105D002AA10FF8002155F7FFC2000080417555FFAA80",
INIT_21 => X"C21EF5D7BC21FFFFFBD55EFAAD1554BA00556AA00AAD140145AA8028ABA002EB",
INIT_22 => X"FFDE00F7842AA00002A80155A2AEA8A10080428A10FFAEBFFEF5D0428B45A2FF",
INIT_23 => X"5568A000000175FFF7D155545F7FBC0010FFAA820AAF7D542155F7D1400AAF7F",
INIT_24 => X"0000000000002AB45082A821EF5D557FF45A2AABFEBA082A975555D55400BA00",
INIT_25 => X"000E38F6D4155504AAA2AEAAB6D0024800000000000000000000000000000000",
INIT_26 => X"05D75E8B6D4120851FFEBD5525C74124B8FC71C71EFA28AAF5E8BFFB6D56DA82",
INIT_27 => X"0014041256DEBA487145F78428ABA147FEDA10080E2AAAA555552400417FC200",
INIT_28 => X"155BE8028A82002EB8FC70024BAEAAB6DB4202849042FA00EB8E0516DE3F5C00",
INIT_29 => X"DFD7550428B55A2F1C71C74975C01FFEBF5D25EFA2D555482085F6FA28AAD147",
INIT_2A => X"4016DE3DF450AAF7F1FDE38FF8A2DA101C2A80145B6AEA8A10080E2DA00F7A0B",
INIT_2B => X"E9557D415B400AA00556DA000004175FFE3D15757DE3F5C0038FFAA800BAF7DB",
INIT_2C => X"000000000000000000000000000002AB7D1C24851FF495F7FF55A2A0BFE921C2",
INIT_2D => X"2D568BEFFFD57FE10002AAABEF0051400AAA2AAAABFF08000000000000000000",
INIT_2E => X"5D5142000007BC20105D5568BFF0004175EFA2D54214508042AB455D517DEBAA",
INIT_2F => X"0AAAE975FFAAD1420005504001FFAA8015545F78028AAA557FFFE00082EAAAAA",
INIT_30 => X"10007BFDEAAA2D557555FF8028A00082EAAB45000028ABAFFFBC20AA08043DE0",
INIT_31 => X"A10002ABFE00F7803FF555D002AB55AAD1575450051401EFA2D5421EFAAD5574",
INIT_32 => X"20BAFFAE820BAFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE10552E82155FFAAA8",
INIT_33 => X"FFF45AA843FE005D2A955FF087BC20AA00517DE000804175EFAAD1555EFA2D14",
INIT_34 => X"000000000000000000000000000000000000000000000028BFF5504175FF087B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000080000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"0001100024A0800000440000000000040088322044200C840000011400151800",
INIT_05 => X"A200014C4000000020000000000B8094020000254C8800000514203000108800",
INIT_06 => X"10000600004B0044020868021428004012120005540812540020008600831000",
INIT_07 => X"00086100043224489428100010811100010001A040003124040CAC6000400009",
INIT_08 => X"00160500090A0282A06400100080C300000005BE0488104C8000000100008800",
INIT_09 => X"00000581041110022000000002002100400080046140011008010100008A0400",
INIT_0A => X"800000000000010180060210200008B2022304080800400007C0100240000000",
INIT_0B => X"0004140000800844522800041004000008000080000400000800000D09240000",
INIT_0C => X"0400004000040000400000000000000000004000020000200000000008010100",
INIT_0D => X"4A00008000000260001001280000C400B0002000000000000000440400000000",
INIT_0E => X"0000000840006000000000001001004004000000000000020100000000000000",
INIT_0F => X"0000000000000000002021000000000000002021000000000000046000240000",
INIT_10 => X"0000000000000000002028000000000000002028000000000000020000008000",
INIT_11 => X"0200000080000000000000000000020001008000000000000000000004000012",
INIT_12 => X"0020000880000000006000400080C0000000000D081202800000000000000000",
INIT_13 => X"0000000100402000000000100000040200100000000000000080009000000000",
INIT_14 => X"0000100000003088014000000000000400000088221100000000000401001000",
INIT_15 => X"4000000800000000048407170500000000000000000400000200000000000000",
INIT_16 => X"00000000023000000220000048240404A010040000008000000000000000020C",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0020014000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000020000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFC0000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"555003DE10A2FBC0000000000000000000000000000000000000000000000200",
INIT_1E => X"BA00003DF555555574AAAAAEAAB45082EBFE000004020AA552E80000F7FBC214",
INIT_1F => X"A00AAFBFDEBA555568BEFA2FBE8A10F7802AA0055003FE10007BE8BEFA2D568A",
INIT_20 => X"55EFF78428BEFAAD17DF55AAAEAAB55552E821FFFFD5555EF552ABDFEF007FE8",
INIT_21 => X"28AAA007FE8A1008002AABA555155400557BC2010557BFFFEFA2FFC20005D2A9",
INIT_22 => X"417555FFAA80155F7843DF455D2AA8B45AAD57FF55A2FBC21FFA28415400FF80",
INIT_23 => X"514200055002AA00AA802AABA002E9740055516AA10FF8002155F7FFC2000080",
INIT_24 => X"00000000000000145AA8028ABA002EBFFFF082EBDEBAA2D1420105D003FFFF08",
INIT_25 => X"412A87010E3F5C0145410E3DE28B6FFC00000000000000000000000000000000",
INIT_26 => X"8147FE8BFFB6D56DA82000E38F6D4155504AAA2AEAAB6D0024B8E381C0A00092",
INIT_27 => X"C74124B8FC71C71EFA28AAF5F8EAA495F68BFFA2F1EFA38E38428A005D0038E2",
INIT_28 => X"FFFBEF5C0000492A955FFF78428BEFB6DB7DF45AAAEA8B6D4120851FFEBD5525",
INIT_29 => X"21EFAA8E10400E38E28ABA147FEDA10080E2AAAA555552400417FC20005D75F8",
INIT_2A => X"0516DE3F5C000014041256DEBA487145F7843FF7D4120A8B6DAAD17FF55B6F5C",
INIT_2B => X"B4202849043FFC7005F4501041002FA38A2842AA82142095428415F6FA00EB8E",
INIT_2C => X"0000000000000000000000000000007155BE8028A82002EB8FC70024BAEAAB6D",
INIT_2D => X"8002AAAA5D2A82000082E95400A2D542155002ABDEBAF7FBC000000000000000",
INIT_2E => X"A2802AA105D002AABA5D7BE8BEFFFD57FE10002AAABEF0051400AAA2AAAABFF0",
INIT_2F => X"F0004175EFA2D54214508042AB455D517DEBAA2D56AABA087BEABEFAAD57DEAA",
INIT_30 => X"00007BC20105D556ABFFF7D142010082A955EFFF8428BFFFFFBFDF55A2AEA8BF",
INIT_31 => X"BEFA2D57DF45F7D1401FFA2AA82000AAAAA8AAA557FFFE00082EAAAAA5D51420",
INIT_32 => X"54AA007BFDE00AAAE975FFAAD1420005504001FFAA8015545F7803FFEF08002A",
INIT_33 => X"AAB45000028ABAFFFBC20AA08043FF55087BD740000043DEAAA2842AA005D001",
INIT_34 => X"000000000000000000000000000000000000000000000017555FF8028A00082E",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000003000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"010108A802BB00080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"8BFA58800005C40A46240252145148B38248030356415A4E62B6FC660F287240",
INIT_05 => X"0F05EA11E570000D610000000710296E542B6E3A825C15FB30A643695BFC2D56",
INIT_06 => X"00000200021100C87570B08224C8AB52C0A8030140BCC0460050690A95C8383D",
INIT_07 => X"76F500240510A00205F0A407D0021A155378900002A002433A0AA00EE6E79564",
INIT_08 => X"00015995440C8327241440096A2800002828123D542910380004E03103624040",
INIT_09 => X"0010222D90409A05B2CB2CA400200209E5601044A24000000462A60018880100",
INIT_0A => X"300000000000259200140001A15000017F0051D0F837248C005514AC40C08205",
INIT_0B => X"395012004240014891801000495D40192D100000000005452D54000C09070003",
INIT_0C => X"6110001100011000110001100011000110001080008800080005202280801080",
INIT_0D => X"BB4000140A80A5C8000102ED0044008004AD324000000008003561180063DB4F",
INIT_0E => X"1400404912AA28AA890BA00000024800480000000000000200802151025062C0",
INIT_0F => X"6D0031F554E11C596A64003195933741477264003195555B418687E358360208",
INIT_10 => X"41CD50A499CF47DCB264003195933741597264003195555B4198843940076D29",
INIT_11 => X"043D400758486A556489347FE5F409CBC1362510695B6288743123C952518520",
INIT_12 => X"B1C74424EAE2992046EB70026486035600CEC45CBCA809654B48163CCC895E1E",
INIT_13 => X"C383298E3A242DEA151848302BFD6D522B10C7EC71F6C1DB071D1216E078C4C1",
INIT_14 => X"8B93D037DAAABC982BE22267A2E2E4F44AA1DC5E37400C9EE1B7B638E8849D23",
INIT_15 => X"86E6A2EE015998B28654565A003F0068E35352C1CAE48BFBF3A6C9B7B286B4DA",
INIT_16 => X"00000000009000040A8000452110A8442040D655602A102A0027E2C423202840",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"B020000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"28A28A28A28F4EF2FC3C34F3CF3C2AC31DF7A22A898D21B4C9838D30B6A7B451",
INIT_1B => X"F4FA3D3E8F4FA3D3E8F4FA68A68A68A68A68A68A68A68A68A68A68A68A68A28A",
INIT_1C => X"FFC00003E9F4FA7D3E9F47A3D1E8F47A3D1E8F47A3D3E9F4FA7D3E9F4FA7D3E9",
INIT_1D => X"AFF80001FF002A80000000000000000000000000000000000000000000000200",
INIT_1E => X"AA552E80000F7FBC214555003DE10A2FBC21FFFFFBFDF45A2D56AB45FFFFD54B",
INIT_1F => X"B45082E974BA5D7BFDF55A2FFFFE005D7BC0010002E954AA087FFFE000004020",
INIT_20 => X"7410FFD1555550000020BAAAFFE8BEFA2D568ABA00003DF555555574AAAAAEAA",
INIT_21 => X"BDEBA555568BEFA2FBE8A10F7802AA0055003FE10007BC0000082A9740055001",
INIT_22 => X"ABDFEF007FE8A00AAFBD55EFAAFBD74105504021FF5D2EAAABAFFFBD55FF002A",
INIT_23 => X"517DF45AAFFFFEAAFFAABFE10007FC00AA087FEAB55552E821FFFFD5555EF552",
INIT_24 => X"0000000000003FFEFA2FFC20005D2A955EFF78428BEFAAD17DF55AAAE820AA5D",
INIT_25 => X"AADB6FB6DFFFBD54AAE38E021FF0824800000000000000000000000000000000",
INIT_26 => X"A1C7FF8E381C0A00092412A87010E3F5C0145410E3DE28B6FFC21C7E3F1F8F55",
INIT_27 => X"6D4155504AAA2AEAAB6D002492482497BFDF45AAFFF8E385D7BC5000002E904B",
INIT_28 => X"010142E90428490015400FFDB555450804070BABEF5E8BFFB6D56DA82000E38F",
INIT_29 => X"DAAAFFF1D55FF002EB8EAA495F68BFFA2F1EFA38E38428A005D0038E28147FC2",
INIT_2A => X"851FFEBD5525C74124B8FC71C71EFA28AAF5D25D7B6F1D54384904021FF5D2AA",
INIT_2B => X"B7DF45AAAE820925D5B7DF45A2F1FDEAAEBAABDE001471C20921475E8B6D4120",
INIT_2C => X"0000000000000000000000000000038FFFBEF5C0000492A955FFF78428BEFB6D",
INIT_2D => X"7FBC2145AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF00000000000000000000",
INIT_2E => X"557FD7410082A800AA557BEAAAA5D2A82000082E95400A2D542155002ABDEBAF",
INIT_2F => X"FFFD57FE10002AAABEF0051400AAA2AAAABFF080000000087BFDF55A2FFE8AAA",
INIT_30 => X"105D002AABA5D7BC20005D2E800BA080417400F7FBD75450800174AAFFD168BE",
INIT_31 => X"4AA0800001EF5D2ABDEBAF7D1575EF082EAAABA087BEABEFAAD57DEAAA2802AA",
INIT_32 => X"0000555568BFF0004175EFA2D54214508042AB455D517DEBAA2D540155F7D155",
INIT_33 => X"955EFFF8428BFFFFFBFDF55A2AE82010557FFDF55A2D57FEAAAAAEBFE1055514",
INIT_34 => X"00000000000000000000000000000000000000000000002ABFFF7D142010082A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000001000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"294ADB4AFFCBF0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"DB7A40806FE4040840EBC563A0150A0926146FECB04196482236FC2005282AE1",
INIT_05 => X"0403DA0383200831C68206D7E6D0250834336D1E81500FDB306045255BFC2076",
INIT_06 => X"D0002200022D1C59E53558D3EBFC6701CBC303163670497AFF00291B3C0E2015",
INIT_07 => X"F81684248A38B022475DCA9BD00116E33CC3821774BB55F53BB42329AA3C0CEA",
INIT_08 => X"1660700CE0641527241060AD844E1C0088001223022D189A2800542219204903",
INIT_09 => X"B6D94C1C1C51DFF881861CBE0305A12A0321810217C01D34EDC98FFA1C8E0000",
INIT_0A => X"F1F1FD8F8FBDE40E001E000B3A5DAADAFDDA5DA79350DF70027CE86F047BEF19",
INIT_0B => X"2DD8141817C00319F8E853E64D73A08BFF00E9A7415606747E6610052CDEE97F",
INIT_0C => X"4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A7800617112E46F05D0",
INIT_0D => X"BFF252D4CFEB69FF7A5F5AFFCCA787F7FE67C2180000006CE8A3F06ABD73DBCF",
INIT_0E => X"94BB02C9F99FD0678B87A0003000D8D02E00000000000000040025D3C21463D6",
INIT_0F => X"6D2BF232221ABD9CA854DFDD64A67D42C0F054DFDD64667D42C063E57A8F7B45",
INIT_10 => X"EFBB5AEDAA504801F054DFDD64A67D42C0F054DFDD64667D42C07237DFE5865F",
INIT_11 => X"3A33DFE58EAE7F5AB50D0806A9A2E0DFFF47DEDC496DA3181A0CC71440F9FBC3",
INIT_12 => X"7056E9C9C3FC95949AEFF556EF9C75E7DCF1EB1B6E6FCDC87CB35FC94B36AECF",
INIT_13 => X"92B29382AF5B6AAAE594A4C0DBFDAD94AA669809809FEFAF4157ADB55572CA52",
INIT_14 => X"BEBF41AE33F32ADD543430808BABAF50E1A5EB4BAEA45A250202FE0ADD39387F",
INIT_15 => X"E83FB669523E865D4B1293AB6B90BF2F0E30EDEFAFD0B3FBD72E9E90D20A003F",
INIT_16 => X"0000000002F840000BCE0B6F67B3F845E017C833F6AAC02B002A2EFF22D4073D",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"CC0C006000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"34D34D34D352324C3434C0EBAEBA21BBE5F04006013DB9880A5D25C3230B88A7",
INIT_1B => X"1A0D06A351A0D06A351A0D34D75D34D34D75D34D75D34D34D75D34D75D34D34D",
INIT_1C => X"FFC00002351A8D46A351A8D46A351A8D46A351A8D468341A0D068341A0D06834",
INIT_1D => X"0007BEAB55FFAA800000000000000000000000000000000000000000000003FF",
INIT_1E => X"45A2D56AB45FFFFD54BAFF80001FF002A821FFFFFFFFFFFFFFBFDFEFAAD14201",
INIT_1F => X"E10A2FBEAB45A28000010082A975EFA2D140145007BC21FF5D2A821FFFFFBFDF",
INIT_20 => X"54AA0855575FFAAD57FE005D7BFFE000004020AA552E80000F7FBC214555003D",
INIT_21 => X"974BA5D7BFDF55A2FFFFE005D7BC0010002E954AA087FD7400082E954AA08001",
INIT_22 => X"5574AAAAAEAAB45082EBFFFFF7D16AB45FFFFEABEF007BD74005555555EFF7AE",
INIT_23 => X"84154BA082E801FFAAFBC0155555568B45552EA8BEFA2D568ABA00003DF55555",
INIT_24 => X"00000000000000000082A97400550017410FFD1555550000020BAAAFFC0145AA",
INIT_25 => X"F7F1FAFD7A2D5400001C7BEDB7DEBA4800000000000000000000000000000000",
INIT_26 => X"F4124821C7E3F1F8F55AADB6FB6DFFFBD54AAE38E021FF0824851FFFFFFFFFEF",
INIT_27 => X"10E3F5C0145410E3DE28B6FFEFB45AA8E070281C20925FFBEDB451451C7BC01E",
INIT_28 => X"4280024924AA1404174AA0055505EFBEDB7AE385D7FF8E381C0A00092412A870",
INIT_29 => X"54005D5B575EFEBAE92482497BFDF45AAFFF8E385D7BC5000002E904BA1C7FD5",
INIT_2A => X"6DA82000E38F6D4155504AAA2AEAAB6D0024BFFD7FFDB6AB7DFFF5EDBC71C7BD",
INIT_2B => X"4070BABEF5C516DAA8A124921C20801FFB6F5C0145555B68B7D4124A8BFFB6D5",
INIT_2C => X"0000000000000000000000000000002010142E90428490015400FFDB55545080",
INIT_2D => X"000155FFF7FBFDFEFFFD568B45AAD5400005D7BFFFEFAA800000000000000000",
INIT_2E => X"FFFFD5545557BC21FF080002145AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF0",
INIT_2F => X"A5D2A82000082E95400A2D542155002ABDEBAF7FBFDF55A2AA974AA5D04001EF",
INIT_30 => X"10082A800AA557BD74BA0004000AA5500174AA0855421FFFFFBEAAAA5D7BEAAA",
INIT_31 => X"BFFF7D57FF455D7FD54105D7BD75FFAAAA80000087BFDF55A2FFE8AAA557FD74",
INIT_32 => X"8BEF000028BEFFFD57FE10002AAABEF0051400AAA2AAAABFF08003FF55F7FFEA",
INIT_33 => X"17400F7FBD75450800174AAFFD1555FFA2AA800105504001EFFFD140145557BE",
INIT_34 => X"0000000000000000000000000000000000000000000000020005D2E800BA0804",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000033FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"0405D434003F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"50805AC31007D6125724029216554A9847669903D640EC8E2001002604503004",
INIT_05 => X"07008000E0EA11803850C800010022660C1C0065003C0404002646DC20A02D40",
INIT_06 => X"30A03A0A138900001127A09234C81FF040000000002C44D620F0228454C83810",
INIT_07 => X"405584280B10014003A8067400920810FF3C72024300A0030048221ACEE383E4",
INIT_08 => X"1000C983E6041505253500F66E620428000B1804000152E52801A20200840900",
INIT_09 => X"0820500B90419005B0C309402030060860E01004A828408800440405E3502940",
INIT_0A => X"A2020010100007865421432121804021C20452880C2D200000045C18C0E0000A",
INIT_0B => X"371097006026226495446E2110AE4417411204400000306B8186185C42900693",
INIT_0C => X"A00308003080030800308003080030800308001840018400400602A018809800",
INIT_0D => X"4008081010108003C000210020460801001FB3650C50DB13111C0D95C20C2030",
INIT_0E => X"14804032007E281F840C00284A17210001060D8306C18360C1380A0260CB9808",
INIT_0F => X"1555D5D79BBEF8E50B041029075982BF3873041029079982BF39748AA0AC8000",
INIT_10 => X"5156AEA479BFD7F7F3041029075982BF3E73041029079982BF3F632C5F96D3C1",
INIT_11 => X"932C5F96A595405FC7F1CFEBC7586C4100A53162B47FD7E39FFEECE159870234",
INIT_12 => X"39464006FE037ACFB88083A99E06271BB0CA207DFDD5920057E0B001B0EBCC79",
INIT_13 => X"6F5DF5CA2A002DD51B6F7FC4A411D1E8D44517F14EAFE36E55150016EA8DB73E",
INIT_14 => X"9DB84953C30351452A13D55CFFA76E928E3891F148B30399F5FB7F28C800DFA0",
INIT_15 => X"110155AC57DFEAEF1005475F1D1F608819CF0EE76E12C824ADD9089715F25FAF",
INIT_16 => X"0D8360D834041A41A0000010180C02801680460FC900052FA10DC0006DA4881C",
INIT_17 => X"D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D836",
INIT_18 => X"8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360",
INIT_19 => X"B000000000000000000000000020D8360D8360D8360D8360D8360D8360D8360D",
INIT_1A => X"1451451451448982C8A82E0820825942495377D9D701DC2E784601F8D187BEF8",
INIT_1B => X"4A2512A954AA5528944A25555145145145555555145145145555555145145145",
INIT_1C => X"FFC00000944A25128944A25128944A25128944A25128944A25128944A2512894",
INIT_1D => X"A5D2E820BA550000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFBFDFEFAAD142010007BEAB55FFAA821FFFFFFFFFFFFFFFFFFFFF7FBD74A",
INIT_1F => X"1FF002A821FFFFFFFFFEFF7D16AB55A2D542000A2D5400BA0800021FFFFFFFFF",
INIT_20 => X"DFFFFFFFC0010F7842AA10F780021FFFFFBFDF45A2D56AB45FFFFD54BAFF8000",
INIT_21 => X"6AB45A28000010082A975EFA2D140145007BC21FF5D2AAABFFF7D168B45AAD57",
INIT_22 => X"BC214555003DE10A2FBEAA00000002010552E95410AAFBD75FF5D7FEAB550051",
INIT_23 => X"04174AA5D00020BA555542145A284155FF5D517FE000004020AA552E80000F7F",
INIT_24 => X"00000000000017400082E954AA0800154AA0855575FFAAD57FE005D7BD740008",
INIT_25 => X"FFFFFDFEFF7FFD74AA552A820AA490A000000000000000000000000000000000",
INIT_26 => X"A080A051FFFFFFFFFEFF7F1FAFD7A2D5400001C7BEDB7DEBA4871FFFFFFFFFFF",
INIT_27 => X"6DFFFBD54AAE38E021FF0824821FFF7F1F8FC7EBD568B7DB6DF47000AADF400A",
INIT_28 => X"BC7E3D56AB7DB6DF78FD7EBF1C2000F78A2DA38E38A021C7E3F1F8F55AADB6FB",
INIT_29 => X"25EF497FEAB7D145B6FB45AA8E070281C20925FFBEDB451451C7BC01EF4124AD",
INIT_2A => X"00092412A87010E3F5C0145410E3DE28B6FFE8A101C0E05010412495428AAF1D",
INIT_2B => X"B7AE385D7FD74381400124825D0A000BA555F47145BE8A105EF555178E381C0A",
INIT_2C => X"00000000000000000000000000000154280024924AA1404174AA0055505EFBED",
INIT_2D => X"A80155FFFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA082A8000000000000000",
INIT_2E => X"F7FBD5410AAFBC00AA002A955FFF7FBFDFEFFFD568B45AAD5400005D7BFFFEFA",
INIT_2F => X"5AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF0000021EFF7D16AB55A2D56ABEF",
INIT_30 => X"45557BC21FF08003FF55AAD168BFFF7FFEAB45AAD140010F7AABFEBAAAAA8214",
INIT_31 => X"4100000154AAA2D1421FF007BE8BFF557BFDF55A2AA974AA5D04001EFFFFFD55",
INIT_32 => X"01EF55516AAAA5D2A82000082E95400A2D542155002ABDEBAF7FBE8A00552E95",
INIT_33 => X"174AA0855421FFFFFBEAAAA5D7BD74BA5D0002010552E820AA5D7BD7545F7AA8",
INIT_34 => X"0000000000000000000000000000000000000000000000174BA0004000AA5500",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000001000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000008128000000000000000000000024001620280000000000354200004008",
INIT_04 => X"000058800004C4024024001210001054B1C822009640000E2000002604003000",
INIT_05 => X"07008000E0200000000000000000200604000000001C04000026400000002C40",
INIT_06 => X"000000000000000004C010B35420015040000000002C42010010200004C83810",
INIT_07 => X"06E200201C00A14080082B26208008A009001201014022404402800408408020",
INIT_08 => X"00004180261C81210031000004340000200008105428020568040213003499C0",
INIT_09 => X"0000000990000000B0C308000000000860200160000000000038380000000000",
INIT_0A => X"10000000000005860000000080A0002060204080000000000004540800000000",
INIT_0B => X"00000000000000020001000022000000000000000000178000F8000101259000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000108000EC000000000000000010004B200000000000000000000000000",
INIT_0E => X"2000000000062801800400000000000000000000000000000000000000000000",
INIT_0F => X"828008084451B81A70AB3006BA0011400760AB3006BA0011400680F020968348",
INIT_10 => X"30B8011204082248A0AB3006BA0011400160AB3006BA0011400084C780687DBA",
INIT_11 => X"64C78068796E80A00802301BC0A7531EDD98E73B02800804620D030F873EB49F",
INIT_12 => X"B0A936B00000002044F091A860700FF9198AA115D5DA37F7A80C8A3604001C06",
INIT_13 => X"0000098551AC9000000000314E01F9F30198600631448410A2A8D64800000081",
INIT_14 => X"1046B2E00303842281C80A23004411AD661891F15148A4420804241526D60000",
INIT_15 => X"66A4A9D335F3D282000C6C5456C84850F61050C411AD6284FDA861682805A04A",
INIT_16 => X"0000000000000000000000000000000000004600C00138000030880042023043",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"9000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C30C30C30C3451046260A9A69A603924554117747E18E0218CC01400163A20C",
INIT_1B => X"26934984C26130984C26130C30C30C34D30C30C30C30C34D30C30C30C30C30C3",
INIT_1C => X"FFC000004C26130984C26130984C26130984C26130984C26130984C26130984C",
INIT_1D => X"A5D2A800105D2E80000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFF7FBD74AA5D2E820BA55003DFFFFFFFFFFFFFFFFFFFFFFFFFD54A",
INIT_1F => X"B55FFAABDFFFFFFFFFFFFFFFFFDFEFF7FFD54BA5D2EA8BFFFF84021FFFFFFFFF",
INIT_20 => X"8B55A2D540010007BEAABAA2AE821FFFFFFFFFFFFFFBFDFEFAAD142010007BEA",
INIT_21 => X"021FFFFFFFFFEFF7D16AB55A2D542000A2D5400BA08003DFFFFFFFFFFFFF7FBE",
INIT_22 => X"FD54BAFF80001FF002ABDFFFFFFFFDFEFA2D56AB45AAFBD74AAFFD5420100804",
INIT_23 => X"FBE8B45AAD568BFFF7FBD74BAFF802ABFFFFAE821FFFFFBFDF45A2D56AB45FFF",
INIT_24 => X"0000000000002ABFFF7D168B45AAD57DFFFFFFFC0010F7842AA10F780155FFF7",
INIT_25 => X"FFFFFFFFFFFFBD54AA5D2A80000412A800000000000000000000000000000000",
INIT_26 => X"7E384071FFFFFFFFFFFFFFFFDFEFF7FFD74AA552A820AA490A38FFFFFFFFFFFF",
INIT_27 => X"D7A2D5400001C7BEDB7DEBA4BAFFFFFFFFFFFFF7FBFDFD7EBF1D24AA5D2AADBD",
INIT_28 => X"FFFFFFBFDFC7E3F5EAB45AAD140000007FEFA92A2AA851FFFFFFFFFEFF7F1FAF",
INIT_29 => X"74AAE3DF400000004021FFF7F1F8FC7EBD568B7DB6DF47000AADF400AA080A3F",
INIT_2A => X"F8F55AADB6FB6DFFFBD54AAE38E021FF0824BDFEFE3F1F8FD7AAD16DB7DBEFBD",
INIT_2B => X"A2DA38E38A125C7E3F1EAB55B6DB6FBD7E3F5D04AAFF8A2DBD7E3A0821C7E3F1",
INIT_2C => X"000000000000000000000000000002DBC7E3D56AB7DB6DF78FD7EBF1C2000F78",
INIT_2D => X"82AA8BFFFFFFFFFFFFFFFFFFFFF7FBD54BA552A80010002A8000000000000000",
INIT_2E => X"A2D5400AA552ABDF55A280155FFFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA0",
INIT_2F => X"FF7FBFDFEFFFD568B45AAD5400005D7BFFFEFAA8028BFFFFFFFDFEFF7FFFFF55",
INIT_30 => X"10AAFBC00AA002ABDFEFF7FBFDF55AAD16AB55AAD140010007BFFE10AAAA955F",
INIT_31 => X"B45A2D57DFFFFFFFD54AAA2FBC20100800021EFF7D16AB55A2D56ABEFF7FBD54",
INIT_32 => X"FF45AA8002145AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF00003FFEFA2D56A",
INIT_33 => X"EAB45AAD140010F7AABFEBAAAAA82155AAD568B55FFFFFDF55A2D1400AAF7AAB",
INIT_34 => X"00000000000000000000000000000000000000000000003FF55AAD168BFFF7FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000002000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"000079800014CC02C034001600000000000000101EC0012EE0C0026E1E80F000",
INIT_05 => X"1F0FF433EFF0440C3902100002203F2EFC040388137C3E20C8EEC00284033CC0",
INIT_06 => X"7000660016490201700000000002FF57C8E8840155FDC0000010E40087D8787A",
INIT_07 => X"4000040007700000000000000001080FF900160000000200C00080001840BFE4",
INIT_08 => X"0009FFBFE5181606000410A4000004202AA8043E0000000000000001209244C0",
INIT_09 => X"0001227FB0000000F7DF78020004011FEFE00000000020031502000083880200",
INIT_0A => X"00000000000015BE0000004000000100000100506002008C2007D5FC80000024",
INIT_0B => X"0020000000000000000000000000000000210018800000000000000010000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000020",
INIT_0D => X"0008000000100000010000002000080101FFB600000000000000000000000000",
INIT_0E => X"0000003007FE29FF800C00000001002040000000000000020480002E42429C00",
INIT_0F => X"000000004D4E180010040000400000001E60040000400000001E6010003C0000",
INIT_10 => X"04000000000094B1E0040000400000001E60040000400000001E608040000004",
INIT_11 => X"0080400002000000000033628000100100000004000000006170C00080010000",
INIT_12 => X"B0020000000000295810000000A100020614148002000000000004307CC3CC00",
INIT_13 => X"000525802000000000014AC000120200000000003F0D800020100000000000A4",
INIT_14 => X"000020020C0C00000000002E2D000001006204040000000005786C0040000000",
INIT_15 => X"004000100A0C0939BEE1810080200000E0CE0EC000010020000000000000AE8A",
INIT_16 => X"000002008040400400C08080000000000049F6FFC01000000000000080080080",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"6902001000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"186186186190324C1090D0F3CF3CD039A060000600704000201120AB02090082",
INIT_1B => X"0C86432190C86432190C86596596596596596596596596596596596596596186",
INIT_1C => X"FFC00002190C86432190C86432190C86432190C86432190C86432190C8643219",
INIT_1D => X"A552A82010080400000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD54AA5D2A800105D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"0BA5500001FFFFFFFFFFFFFFFFFFFFFFFBD54BA552A8001000003DFFFFFFFFFF",
INIT_20 => X"FFEFF7FFD74BA552E801FF002E821FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E82",
INIT_21 => X"BDFFFFFFFFFFFFFFFFFDFEFF7FFD54BA5D2EA8BFFFF843FFFFFFFFFFFFFFFFFF",
INIT_22 => X"142010007BEAB55FFAA801FFFFFFFFFFFFFFBFDFEFFFD542000082EAAB55AAAA",
INIT_23 => X"FFFFFFFF7FBFDF55AAD140000087BE8B55F784021FFFFFFFFFFFFFFBFDFEFAAD",
INIT_24 => X"0000000000003DFFFFFFFFFFFFF7FBE8B55A2D540010007BEAABAA2AE975FFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA552A820001400000000000000000000000000000000000",
INIT_26 => X"81C0038FFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2A80000412ABFFFFFFFFFFFFF",
INIT_27 => X"EFF7FFD74AA552A820AA490A021FFFFFFFFFFFFFFFFFFEFF7FBD74BA5D2A8002",
INIT_28 => X"FFFFFFFFFFFFFFFBFDFEFFFFFD54BA5D2A801C7142E871FFFFFFFFFFFFFFFFDF",
INIT_29 => X"0010142AAFB7DBEAEBAFFFFFFFFFFFFF7FBFDFD7EBF1D24AA5D2AADBD7E38438",
INIT_2A => X"FFFEFF7F1FAFD7A2D5400001C7BEDB7DEBA4871FFFFFFFFFEFF7FBF8FD7E3D14",
INIT_2B => X"FEFA92A2AA925FFFFFFFDFEFE3F1FAF45A2D142010087FEDB55F78A051FFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFBFDFC7E3F5EAB45AAD140000007",
INIT_2D => X"02ABFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005D040000000000000000",
INIT_2E => X"F7FFD74AA5D2A800BA550428BFFFFFFFFFFFFFFFFFFFFF7FBD54BA552A800100",
INIT_2F => X"FFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA082A821FFFFFFFFFFFFFFBFDFEF",
INIT_30 => X"AA552ABDF55A2802ABFFFFFFFFFEFF7FBFFFFFF7FBD74BA552A80145552E955F",
INIT_31 => X"FEFF7FFEAB45AAD1420105D2ABFFFFFFAEA8BFFFFFFFDFEFF7FFFFF55A2D5400",
INIT_32 => X"DF55F7AE955FFF7FBFDFEFFFD568B45AAD5400005D7BFFFEFAA80175FFFFFBFD",
INIT_33 => X"6AB55AAD140010007BFFE10AAAA821EFF7FBFDFFFAAD168B55A2D542010007BF",
INIT_34 => X"00000000000000000000000000000000000000000000003DFEFF7FBFDF55AAD1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"084A76341244919000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"000079800014CC03C075161E001118653D2408041FC004AEF000816E1C11F541",
INIT_05 => X"3F0F807BFFE000240100004683103E7FFE02482553FC3C0204EFC25010143CC0",
INIT_06 => X"1100441004201014B1709C910102FF5FC0A0000101FFE4036450E08247F87870",
INIT_07 => X"08750504800680102542AD800504530FF9061E8026998E9A00402CC25BD0FFFC",
INIT_08 => X"0011FBFFE04691A5A00101818A6800088228000001A044C8168480D010F200AA",
INIT_09 => X"B6E85A7FF080AC70FFDF78220010841EFFE7116E144071268DFD3E4C24040100",
INIT_0A => X"3151518A8A31B7FE00040009814C089202225412115428C03BC7D7FC15025B1A",
INIT_0B => X"1B1883007104032901CC63410ABD249C4B338934404037FC8BFE18008083B444",
INIT_0C => X"D9228D9228D9228D9228D9228D9228D9228D99146C9146C84006309044081A00",
INIT_0D => X"48000201800500941044312000900D4621FFBE00080081529904595123203040",
INIT_0E => X"308162029FFEADFF8050250010030165290008800440022201082401A002000C",
INIT_0F => X"5001318048A004A6C0D2820302C005A83480D1820302A009B02B101390C0CB28",
INIT_10 => X"485101408904831400D1820302C005A83480D2820302A009B02B021A85C09411",
INIT_11 => X"FA1A85C08834600024D052C1051E0B92D400360520202682C19024B6164E3004",
INIT_12 => X"C1B0D6404093E22A2012418A9D1D44ADD9E0F174103820101C0B8160D5516259",
INIT_13 => X"6C88660D8AA288209E615100280DA0052000C5006402000206C55144104D510C",
INIT_14 => X"024500A0D50020C04023033C52009144231D902818100C90058010361AC80812",
INIT_15 => X"198A12202386454988140600C0181500A13E830011008B0374007000B4E0CD00",
INIT_16 => X"008020080224004002000000703804008001F7FFF01B982B01258088C008CC41",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"F000000000000000000000000020080200802008020080200802008020080200",
INIT_1A => X"7DF7DF7DF7DFFFFEFEFFFE79E79FFFF3BC1FF3FDDFEFFFBEFFE7DF84081EFEFB",
INIT_1B => X"FEFF7FBFDFEFF7FBFDFEFF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF",
INIT_1C => X"FFC00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"A5D2E80010000400000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA552A8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"0105D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E80010552EBFFFFFFFFFFF",
INIT_20 => X"FFFFFFFBD54BA5D2E82010002ABDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A80",
INIT_21 => X"001FFFFFFFFFFFFFFFFFFFFFFFBD54BA552A800100000001FFFFFFFFFFFFFFFF",
INIT_22 => X"BD74AA5D2E820BA5500001FFFFFFFFFFFFFFFFFFFFF7FBD74BA5D2E800BA5D00",
INIT_23 => X"FFFFFFFFFFFFFFEFF7FBD74AA552A800BA5D2E821FFFFFFFFFFFFFFFFFFFFF7F",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFEFF7FFD74BA552E801FF002E975FFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E800000800000000000000000000000000000000000",
INIT_26 => X"05D2ABFFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8200014003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFBD54AA5D2A80000412ABDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2E8000",
INIT_28 => X"1FFFFFFFFFFFFFFFFFFFFF7FBD54BA552E82028002AB8FFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74AA5D2E800AA5500021FFFFFFFFFFFFFFFFFFEFF7FBD74BA5D2A800281C0000",
INIT_2A => X"FFFFFFFFFFDFEFF7FFD74AA552A820AA490A071FFFFFFFFFFFFFFFFFFEFF7FBD",
INIT_2B => X"A801C7142E955FFFFFFFFFFFFFFFFDFEFF7FFD54BA5D2E80082492E871FFFFFF",
INIT_2C => X"0000000000000000000000000000038FFFFFFFFFFFFFFFBFDFEFFFFFD54BA5D2",
INIT_2D => X"D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008000000000000000000",
INIT_2E => X"FFFBD54AA5D2E800005D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF7FBD54BA552A80010002ABDFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"AA5D2A800BA5504021FFFFFFFFFFFFFFFFDFEFF7FBD74AA552E820BA002AA8BF",
INIT_31 => X"FFFFFFBFDFEFFFFFD54BA552E800BA5D04021FFFFFFFFFFFFFFBFDFEFF7FFD74",
INIT_32 => X"0000082A955FFFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA082A955FFFFFFFF",
INIT_33 => X"FFFFFF7FBD74BA552A80145552E975FFFFFFFFFEFF7FBFDFFFFFFBD74AA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000002ABFFFFFFFFFEFF7FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"431965109E4481D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"492C0020220001010E4916C884DCD607E5EC2A344103E48003D0800023D0072C",
INIT_05 => X"00107C441001100D620A06D683018001023D37E5088043620101179092540112",
INIT_06 => X"401002010042384D223C19C3552800081ADA0E054402365774611E047020008E",
INIT_07 => X"491EC04ED017AB5497EB923F08182E20020689B735011FBFE7BC062602944019",
INIT_08 => X"154A00401D4425ADA9035BE19C8F9442A8801200F4C9D7AC8093A051727B2AC3",
INIT_09 => X"9A50020040E48D50080002B00A0C00801014541E9504703680017F6CB4050700",
INIT_0A => X"8151538A8A738041C23020131A80CFDFF3FE509A907C6AC05040220409009031",
INIT_0B => X"2D040050110081E9528963546278008AA80381B4000500026800000109379864",
INIT_0C => X"1C2A81C2A81C2A81C2A81C2A81C2A81C2A81C9540E1540E00140000610000320",
INIT_0D => X"594A06870A9CA0D458D131652A154D46B6000850800801628013456520CA0928",
INIT_0E => X"02080448C00044000A1EC1C44140D101A54280A14050A028500A84F02842A24C",
INIT_0F => X"0061338359E0C4E6C256690581800F1C3E82562B0581200F1C3F081456022804",
INIT_10 => X"2C438100AB8581B602562B0581800F1C3E8256690581200F1C3F1238473F1210",
INIT_11 => X"2238473F0E1050083750B3E4275F829547008600C030374361FA2CEE046D4812",
INIT_12 => X"C1128C4CC012A66F61154C019511628756231018500C00203E13806156516078",
INIT_13 => X"54CDE608AA612C0096C37B00D1724801A0009C606D1221D104553096004B61BC",
INIT_14 => X"870B012A41E0F0600035842E7601C2C4AC68A98810080AA825A8902251899802",
INIT_15 => X"58234A89637E00D0A1080301401C390320188321C2C0B13890105800D520AF94",
INIT_16 => X"8822088222F110111B281A54753AA004002601001918008C10912A4440B24E8B",
INIT_17 => X"8220882208822088220882208822088220882208822088220882208822088220",
INIT_18 => X"2008020080200802008020080200802008020080200802008022088220882208",
INIT_19 => X"E82891448000000001FFFFFFFFC8020080200802008020080200802008020080",
INIT_1A => X"3CF3CF3CF3DFFBFEFEBEEEFBEFBEFBEBFDF7F7FBDFD1FE3EFBD7ADFBF7EFBEFB",
INIT_1B => X"FE7F3F9FCFE7F3F9FCFE7F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"FFC00001FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"A5D2E82000000000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8000008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74AA552E8000055003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A82",
INIT_21 => X"BFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E80010552EBFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD54AA5D2A800105D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A82000552A",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD54AA5D2A800005D2EBDFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000000001FFFFFFFFFFFFFFFFFFFFFFFBD54BA5D2E82010002AA8BFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100004000000000000000000000000000000000",
INIT_26 => X"008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA552A8200014003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E800105D043FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"54AA5D2A82010552EBDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2E800005D2ABF",
INIT_2A => X"FFFFFFFFFFFFFFFFFBD54AA5D2A80000412AB8FFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E82028002AA8BFFFFFFFFFFFFFFFFFFFFFFFBD54BA552E80038492EB8FFFFFFF",
INIT_2C => X"00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFF7FBD54BA552",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000040000000000000000",
INIT_2E => X"FFFFD74BA552A8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E800000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005D043FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"AA5D2E800005D2EBDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA552E8001055003FFF",
INIT_31 => X"FFFFFFFFFFFFF7FBD54BA5D2A820105D2ABDFFFFFFFFFFFFFFFFFFFFFFFFBD54",
INIT_32 => X"00AA082EA8BFFFFFFFFFFFFFFFFFFFFF7FBD54BA552A80010002AA8BFFFFFFFF",
INIT_33 => X"FDFEFF7FBD74AA552E820BA002AAABFFFFFFFFFFFFFFFFFFEFF7FBD74BA552E8",
INIT_34 => X"0000000000000000000000000000000000000000000000021FFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"2C4360101A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"00017B810015DC03D034201E14000036486008101FC0002EE006297E1C05F561",
INIT_05 => X"BF0F817FFFE80100004044800080BEFFFC0248005FFC3C18A5FFC2444484BCC0",
INIT_06 => X"B0801408110000109127E0500002FFDFC000000001FFC0832050E00047F97870",
INIT_07 => X"00D1D72040048D00388387D03D0E591FFD201F862691DFBE077C2BC45B40FFE4",
INIT_08 => X"001FFBFFEC440501A5604B31062356282AA84200D12342113EDC400000045828",
INIT_09 => X"25A890FFF0002023FFDF79000000000EFFE309606020008005FC000000402000",
INIT_0A => X"30000000000037FF50010103134CAFDF03BA18000F39A0106F87D7FA84024B02",
INIT_0B => X"1B188300624483890564084198AD249C43300C00415037FC83FE1840C0902400",
INIT_0C => X"C1010C1010C1010C1010C1010C1010C1010C10086080860840063090442A1800",
INIT_0D => X"0001403000100200180480000095280001FFBF040C40C81119A41C1443243050",
INIT_0E => X"32A163821FFEAFFF805025E00853B92588000400020001000020A80180080020",
INIT_0F => X"90401486148484054395E27E428002A4200397E07E422002A420100382FCC308",
INIT_10 => X"641100C0788417000397E07E428002A4200395E27E422002A420110A51C01C05",
INIT_11 => X"C90A51C01A2490040590C08120558C1759BE1C05A0400383808800DA1929F728",
INIT_12 => X"00CE720000136006000215EA0A4833A32C8832050028603050014031B3950000",
INIT_13 => X"6C00C006658280009A2030108B14AC05C00112405222088B8332C140004D1018",
INIT_14 => X"A2659196B6808060201281004228996085F10020180C030880D11019CE400002",
INIT_15 => X"0108152A49DC7143F01C04240030720641E0A028996483A17204680410A04104",
INIT_16 => X"040100401000080080000000000002001201F7FFC0011C2F81A48080CA32800A",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_19 => X"0000000000000000000000000000401004010040100401004010040100401004",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000020000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFC0000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2A8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E80",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8000008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA552A8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A820000004",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA552A8201000043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E8000055003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA552A8200008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001008043F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA552A8200014003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E800105D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E820101C003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552",
INIT_2D => X"0043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA552A8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001008043FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74AA552A8200008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"200055043FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005D043FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD54AA552E8001055003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA552E8",
INIT_34 => X"00000000000000000000000000000000000000000000003DFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"00003A2E200811000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"000079800014CC03C034001E04010850300000101FC0002EE000006E1C00F500",
INIT_05 => X"1F0F8033FFE000000000000000003E2FFC024800137C3C0000EFC00000003CC0",
INIT_06 => X"000000000000000091C115500002FF5FC000000001FFC0000010E00007F87870",
INIT_07 => X"10E600084002040A10812A000500590FF9001F95406A8000037230C01840FFE0",
INIT_08 => X"0001FBFFEC4695A501604A000C7585080002C200408102F16C0184800026C92C",
INIT_09 => X"24A8107FF0000000FFDF78000000000EFFE001600000000005FC000000000000",
INIT_0A => X"30000000000037FF4000000AA0354000019C4000012800002387D7F804024B02",
INIT_0B => X"1218830060040A04000400000801241443300800404037E883FE180000000000",
INIT_0C => X"C1000C1000C1000C1000C1000C1000C1000C1000608006084006301044081800",
INIT_0D => X"00000004800B0000000000000000000001FFBE00080080101904181003003000",
INIT_0E => X"B08062021FFEADFF800020800000002088000000000000000000200180000000",
INIT_0F => X"D0210840009181008024A00043601100210024A00043C0110020901382CCCB28",
INIT_10 => X"0C920180040A03080024A00043601100210024A00043C01100209240C840C201",
INIT_11 => X"1A40C840A604E0080820009908008341B000A821207008200289001006832086",
INIT_12 => X"0166B40600800082041205EC00044C1ACB66C37542082030281E058000101281",
INIT_13 => X"0010480B27A004300004103160DB3005E000618040C022000593D00218000209",
INIT_14 => X"880012BBFF20406040084210C062000C2A2DDD00180C04504086002CD680C010",
INIT_15 => X"4106020804295C98F80400008040CC0582169022000C2876C404780028500160",
INIT_16 => X"000000000000000000000000000000000001F7FFC001B823018F008800088052",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"C800000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"7CF7CF7CF7D933CC3090CABAEBAFF969319815DD5EDCF9822659AE7B095A220C",
INIT_1B => X"1E0F0783C1E0F0783C1E0F7DF7DF7DF3CF3CF3CF3CF3CF7DF7DF7DF7DF7DF7CF",
INIT_1C => X"FFC000003C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C",
INIT_1D => X"A5D2E82010080400000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"00000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E800000800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8001000003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100804000000000000000000000000000000000",
INIT_26 => X"000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"A8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000043FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008040000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8000008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"000008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2A8001008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00002000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"924279824C94CC1BE0B4001F20000000020380401FE0082EF000106E1C00F500",
INIT_05 => X"1F0F8033FFF048202582800100523E2FFE024820137C3C0040EFE02000003CE4",
INIT_06 => X"F10466105670019C900000100002FF5FC0E0801101FFC0000010E08A07FC7870",
INIT_07 => X"0000040000000000000000000500590FF9001F0000000000033020C01840FFFC",
INIT_08 => X"0001FBFFFD0004000100502000011400000282004001020000000001009015C0",
INIT_09 => X"2CB8DA7FF8004000FFDF7C062031863EFFF75D78004001010DFC000020050100",
INIT_0A => X"30000000000037FFC00602000000000001980400002800032387D7FE94FBEF2B",
INIT_0B => X"9258830060040200000400000801243443B00808404037E883FE180C00000000",
INIT_0C => X"C1000C1000C1000C1000C1000C1000C1000C10006080060840077330C4889CC2",
INIT_0D => X"0000000000000000000000000001280001FFBE00080080101904189003003000",
INIT_0E => X"30A063021FFEADFF805025C0304001E58906088304418222C108A009A0904000",
INIT_0F => X"1000000000100100000480000200100000000480000200100000100380F0C308",
INIT_10 => X"0010000000080000000480000200100000000480000200100000000040400000",
INIT_11 => X"0000404000040000000000080800000110000000200000000200000000012000",
INIT_12 => X"00021000000000800002018C0100000208000008001220000000040040000080",
INIT_13 => X"0010000020800000000400000010200200000000008002000010400000000200",
INIT_14 => X"0800000210000080010000008002000000210000201000000002000042000000",
INIT_15 => X"0184000000084000000006050000000002000002000000204000000000000020",
INIT_16 => X"08822288226410410346010000000400A011F7FFE00318230104008000008000",
INIT_17 => X"8822088220882208822088220882208822088220882208822088220882208822",
INIT_18 => X"8220882208822088220882208822088220882208822088220882208822088220",
INIT_19 => X"0404000017FFFFFFFFFFFFFFFFE0882208822088220882208822088220882208",
INIT_1A => X"492082492085048029890AD34D35FDD04A165129432D518B45265EFC30760AED",
INIT_1B => X"C46231188C46231188C462492492492492492492492492082082082082082082",
INIT_1C => X"FFC000058AC562B158AC562B158AC562B158AC562B158AC562B158AC562B158A",
INIT_1D => X"A5D2E820100800000000000000000000000000000000000000000000000003FF",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100000",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000043FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"4A53D958C50000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"DBFAFBD7FB1CDEBEF1BE17F7AC88042787FBFFF8FEE9FF7EE6F4C0EE1FFAF869",
INIT_05 => X"5F0FFEB3EFFEFFBDA7F7FED508707E2EFEBF6FFEB37C3FF302EEEDFF9B487CF6",
INIT_06 => X"74EADE4EBDFDAC9930F6F8129E3FFFF7C3E3A74667FDDB7FB870FF30FFDEF87F",
INIT_07 => X"8173840C07783060C72DF7D828912E6FFB80162776F3BFB7077E82255E40BFEF",
INIT_08 => X"4769FFBFE43C872321367036163F1C0820A3063F460D1AEFC000060042648C41",
INIT_09 => X"BEFB967FBD13D981F7DF7D7E6171AF3FEFE8A3E679FAC1FD1FFFBEB000763A84",
INIT_0A => X"F3A3AD1D1DAD7FBE7D67D7F3BB79CFFB83BF14EC1E7D7300B017F5FFE6FBEF73",
INIT_0B => X"52199F58F6EE6F5E7FAC4C03DB856CD4CF720FE8C4427FF8CFFE38FF7F6BD928",
INIT_0C => X"F78C0D78C0D78C0D78C0D78C0D78C0D78C0D7A606BC606B8C56F7730ECCDBDF1",
INIT_0D => X"EA035CF6100C0E60FB9FC3A80EF69A04DFFFF7FF5E75FF341B867D3683A03A40",
INIT_0E => X"36B867027FFFF9FF8FAFAA3ADEBFB9726BAF5FD7AFEBD7F7EFFD7ACDB7F947F0",
INIT_0F => X"10003E020080A40403E8BD8002000FC02003E8BD8002000FC02010979AFFE36C",
INIT_10 => X"80100000EE00034003E8BD8002000FC02003E8BD8002000FC020037B0040A000",
INIT_11 => X"037B0040C00400003D80008160400FD81341C00020003B80008C00801EF02853",
INIT_12 => X"01F1190981038406809677FA080468C46A81080581002000780C8001C8100201",
INIT_13 => X"7080D00F90D162001C803411FC0024080001F80040026C0807C868B1000E401A",
INIT_14 => X"B02013F810503A00003E020042AC080CEB01228A80000F600080123E23213040",
INIT_15 => X"61F810087520750001064180807868000110C02C080CFA0042400000F8800105",
INIT_16 => X"5FD7F7FDFF7EFEEFF3EEC3FF7FBFFBCB7FFFFEFFE00BFF7FEBF420800EC0CBEE",
INIT_17 => X"FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F",
INIT_18 => X"D7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5",
INIT_19 => X"6DAE443237FFFFFFFFFFFFFFFFF5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5F",
INIT_1A => X"4D34D30C30DD795EAA6AFC38E38EA3AB788962B79E923C2CD990A7D3B4A9FC37",
INIT_1B => X"26130984C26130984C26130C30C30C30C30C30C30C30C30C30C30C30C30C30C3",
INIT_1C => X"FFC000004C26130984C26130984C26130984C26130984C26130984C26130984C",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"0842D85841000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"DBEAE5D6D91C2EBCE1B21EA72C00000007FBE7C8F8E9EF79E6D440E91FDAE061",
INIT_05 => X"5C8FFCB38FF6B68984B5BCE408347E28FEBF6FEEB3723F7102E8EDBF8A4872F6",
INIT_06 => X"946ACF46ACE0841A00006A089E3FFF27C3032646EFF1DB7FA868FE30EF1CE47E",
INIT_07 => X"8000000A20083060C00C81882A008C6FF880060424B39FB6037F00051C003FE0",
INIT_08 => X"4761FA3FE4010440410844060001040A00002200460D1A060000050400000010",
INIT_09 => X"FEEB027E390A4881C7BEFC5F6171CE2F8FE823E778DAC16C1FFBBC9000315895",
INIT_0A => X"F606013030213C3E2D62D6E21259CFDB039E806C024531008017C1F826FFEF41",
INIT_0B => X"5219AB5AF86F7D5E382A440349816DD4C7560B60D4427FF0C7FEBABF3F6BD108",
INIT_0C => X"E3440C3440C3440C3440C3440C3440C3440C3C2061A2061AD46FF730E5CCBCD5",
INIT_0D => X"6203E8FC10080A20ED1D41880CC61A044DFFC6EB5AB5B7941BC63F1683803C00",
INIT_0E => X"B88572023FFE91FF98AEAA1AC6AC9A3A4AAD5B56ADAB56D5AFD572C597B14750",
INIT_0F => X"10003E020000260403C8948002000EC0000BC8948002000EC00010878AC3CB8A",
INIT_10 => X"80100000EE0000400BC8948002000EC0000BC8948002000EC000097B00402000",
INIT_11 => X"017B0040400400003D80000070400DD81041400020003B80000410801AF02041",
INIT_12 => X"05D11101010384008086378A080428C46A80080081002000780C800188000301",
INIT_13 => X"7080102E909042001C800409FC0020080001F80000007C0807484821000E4002",
INIT_14 => X"F02003F810100A00003E020000BC0808EB01020280000F60000002BA22202040",
INIT_15 => X"21F810007520750000024080807868000100403C0808FA0040400000F8800001",
INIT_16 => X"5B56D5B5EF3AF6AF6389C2FE128971AB2DDDF8FFE0031B776BF4208006C0C926",
INIT_17 => X"B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D",
INIT_18 => X"56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5",
INIT_19 => X"238B443A3FFFFFFFFFFFFFFFFFD5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B",
INIT_1A => X"00000000000F0080397908000000A4805F09C42D0200903950C086D420010825",
INIT_1B => X"8040201008040201008040000000000000000000000000000000000000000410",
INIT_1C => X"FFC00005028140A05028140A05028140A05028140A05028140A05028140A0502",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100804",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"461080404900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"00800040110102000902002000888400081045A8A00003C00000500000080008",
INIT_05 => X"0000000000024CA0A0101800032000400000000B800000014000000B08180000",
INIT_06 => X"0020280202802C00020800008A14002011110012220009A88800009A88000000",
INIT_07 => X"8108044200091224484510201000204000800020410000000080000104000009",
INIT_08 => X"132800000140200808021006108010422AAA8000224489028492201140092240",
INIT_09 => X"0001C800004080A0000002480B04008100011000088800081002C19020150B00",
INIT_0A => X"4353529A9A528000040040702080000000400064080011001050000200000018",
INIT_0B => X"01400048012220122A0004168110400004000040811600000400001036584108",
INIT_0C => X"36050160501605016050160501605016050160280B0280B00120008430660210",
INIT_0D => X"2A000C4210040860B188C0A8065302005A0040390010120500002002C0040010",
INIT_0E => X"8221050060001000028000080205001066000100008000400490020402010530",
INIT_0F => X"000000000000A00000081480000001400000081480000001400000800C010820",
INIT_10 => X"8000000000000240000814800000014000000814800000014000000100002000",
INIT_11 => X"000100004000000000000001400000080041400000000000000C000000100041",
INIT_12 => X"000101010100000480802A400000004000000800810000000000000048000000",
INIT_13 => X"0000900010104200000024000400000800000000000244000008082100000012",
INIT_14 => X"1000004000100A00000000000284000040000202800000000000120020202040",
INIT_15 => X"2050000010000000000240800000000000104004000040000040000000000005",
INIT_16 => X"010040108408420430E699AA42A1508104EA08000000810020000000044001AC",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"0506117080000000000000000000100401004010040100401004010040100401",
INIT_1A => X"4104104104006C1A8283AC618618EF10C0422205822140048D2E581E80DEC4D2",
INIT_1B => X"C06030180C06030180C060410410410410410410410410410410410410410410",
INIT_1C => X"FFC0000582C160B0582C160B0582C160B0582C160B0582C160B0582C160B0582",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0401D940CD0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"49B87A417315D20A313E17F1800000058013DDF8BE21F36E02F0D06E03E8F800",
INIT_05 => X"1F007E33E01A4D9C87525E5101603E6E023D27DA937C03E340EE25CB9B483C12",
INIT_06 => X"F0A05A0A15AD0C0130F6F0128A16FFF001E1870223FC3BFC98101F109FC6780F",
INIT_07 => X"8073800407781020476467D008910A4FFB80100332D1AE93059282215E408006",
INIT_08 => X"0221FF80003C832320342036063F08000001063F42050AEB4000221000248C01",
INIT_09 => X"9A51547F8C1111A0F041056A0100A11FE000916249A800B915FE82B020522900",
INIT_0A => X"42A2AD1515AD5780540541619968C76980E914E4163D53002017F405C409A42A",
INIT_0B => X"0140140816A22B126DA40C03531440800C2005C8800217F80C000055FF7C4928",
INIT_0C => X"268D0068D0068D0068D0068D0068D0068D006A68034680300021410028450530",
INIT_0D => X"AA01587410080C60AB0F42A804628200DBFFF13D04505B2500806522C0A40A50",
INIT_0E => X"941922006FFFF8000F8F80281A16A1504302058102C0816244B82A0CA25907D0",
INIT_0F => X"000000000080A40000283D80000001402000283D80000001402010901A7D6944",
INIT_10 => X"800000000000034000283D80000001402000283D80000001402002010000A000",
INIT_11 => X"02010000C000000000000081600002080341C00000000000008C000004100853",
INIT_12 => X"0021090981000006809076B20000404000010805810000000000000048100200",
INIT_13 => X"0000D0011051620000003410040004080000000040026C00008828B10000001A",
INIT_14 => X"B000104000503A000000000042AC00044000228A800000000080120421213040",
INIT_15 => X"607800081000000001064180000000000010C02C000440000240000000000105",
INIT_16 => X"05816258964C4A44A0C689FF3F9FFEC5D6DBFE0020096528A0B000000CC043EC",
INIT_17 => X"5816058160581605816058160581605816058160581605816058160581605816",
INIT_18 => X"8160581605816058160581605816058160581605816058160581605816058160",
INIT_19 => X"F506003017FFFFFFFFFFFFFFFFE0581605816058160581605816058160581605",
INIT_1A => X"5D75D75D75DFFFFEFCFDF7FFFFFF5DE7FC3DF3F2DDCFFFBEFFCF1F84421FFEFF",
INIT_1B => X"EFF7FBFDFEFF7FBFDFEFF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF75D7",
INIT_1C => X"FFC00007DFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDF",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"E800000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"3CF3CF3CF3DD7FDEBAFAFEFBEFBFFBFBB9DFF7FFDFF3FC3EFFF7FDFBBDFFFEFF",
INIT_1B => X"FE7F3F9FCFE7F3F9FCFE7F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"FFC00001FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"08425818000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"DB6A618248140C18E0B016872400000007EBA24058E1ECA8E2D400681FD0E061",
INIT_05 => X"1C0FFC338FF01009048084C400103E28FE3F6FE513703F7000E8E5B4825030F6",
INIT_06 => X"100046000460001800006800142AFF07C202060445F1F2572060FE82671C607E",
INIT_07 => X"00000008800020408008818838000C2FF800060424B39FB6037E000418003FE0",
INIT_08 => X"0441FA3FE4000400010040000001040880000200440912040000040000000000",
INIT_09 => X"BEE8027E38004801C79E7C162231862E8FE00166704041240DF93D0000000000",
INIT_0A => X"B00000000000343E002202021259CFDB039E0008024520000047C1F804FBEF01",
INIT_0B => X"121883107044094C1028400548812494C3120920404437F0C3FE180D89279000",
INIT_0C => X"C1000C1000C1000C1000C1000C1000C1000C18006080060840477330C4889CC0",
INIT_0D => X"400340B400080200481501000884080405FF86400800811019861D1403803800",
INIT_0E => X"308062021FFE81FF880EA000400098200C04080204010200810020C180904240",
INIT_0F => X"10003E020000040403C0800002000E800003C0800002000E8000100780C2C308",
INIT_10 => X"00100000EE00000003C0800002000E800003C0800002000E8000017A00400000",
INIT_11 => X"017A0040000400003D80000020400DD01000000020003B80000000801AE02000",
INIT_12 => X"01D01000000384000006118A080428846A80000000002000780C800180000201",
INIT_13 => X"7080000E808000001C800001F80020000001F8000000280807404000000E4000",
INIT_14 => X"A02003B810000000003E020000280808AB01000000000F600000003A02000000",
INIT_15 => X"01A81000652075000000000080786800010000280808BA0040000000F8800000",
INIT_16 => X"08020080223010010308025410082404A015F0FFE003182701B420800280C802",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_18 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_19 => X"0008004017FFFFFFFFFFFFFFFFC0802008020080200802008020080200802008",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFC0000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"441406267B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"0005802424830120024121209088809DF81454ACA01E03501D0A3B91E00F0A00",
INIT_05 => X"E0F001CC00012034C20B0232838F80D001C0100AEC83C008EF101A034C8CC300",
INIT_06 => X"2F1620F1721BA346AA2C95C5CB1400000161F84322000DA8C40F003C80030780",
INIT_07 => X"5939F36677EE1C387777622717EF711004A6818111086008E080FDC305940018",
INIT_08 => X"13160400195E83A3A0F61BC3929ECB622AABF5FF83860CEB164833F179B48CEE",
INIT_09 => X"01036D8004FDB47600000229410C61010016DC998C84B0128202C0DCB48F05D5",
INIT_0A => X"4400402A0A37000182502440888420247041E876810099D35F900002DB00105C",
INIT_0B => X"AD4434020CA2E0B32B01A752B078412A24818094151348062400E2A034D86444",
INIT_0C => X"3E2781EA781E2781EA781E2781EA781E2781C33C0613C0E21028840239452116",
INIT_0D => X"394818429A95E954868AD0E52273F54258000080808900C3807122C3E04E0338",
INIT_0E => X"8E3B15C94001120055704DC4A1624487E2489024481224091282C4300942A194",
INIT_0F => X"C06101C55D65C3E3F01F52FFC1E0013C1F801F52FFC1E0013C1F8090423D38A1",
INIT_10 => X"ECC381C0118796BE001F567FC1E0013C1F801F567FC1E0013C1F9085DFBF7E15",
INIT_11 => X"F885DFBF7E30F00C0270F3751F1FD00FECBF7E25C0700463E17B2C7F811FD7AD",
INIT_12 => X"C40FE6474190626D6491063597F9177B956EF378D33E4030061341F077C571F8",
INIT_13 => X"0C4DAE207F328E3082636B2807FFD80FE00007E03F7207D3E03F9167184131B5",
INIT_14 => X"1F4FE047EFA0CAE06101C53E3647D3F144FCDD22B81C0098E57D9081FCE8C852",
INIT_15 => X"38574FF31ADF08DBF81846A540049707E0FE3307D3F141FFB45478040570EED4",
INIT_16 => X"90240902C189601208A1102B4AA5584B4068000019A80098120BCA4C617635C9",
INIT_17 => X"0240902409024090240902409024090240902409024090240902409024090240",
INIT_18 => X"2409024090240902409024090240902409024090240902409024090240902409",
INIT_19 => X"9AA09426A8000000000000000009024090240902409024090240902409024090",
INIT_1A => X"104104104104431042720EE38E38AAF9A93E7131C136AD8E9B562CF03B2E8E78",
INIT_1B => X"F87C3E1F0F87C3E1F0F87C104104104104104104104104104104104104104104",
INIT_1C => X"FFC00001F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0",
INIT_1D => X"AAAAABDEBAF7AE8000000000000000000000000000000000000000000000C200",
INIT_1E => X"EFF7D142145A2AE800BA08514214555517DEAA5D7BFFEAAF7803FEBAF7FFD74B",
INIT_1F => X"E00A2FBD75FFFF84001550851555FF55517FE000055421FF00557DF45A2D5401",
INIT_20 => X"74BA552EBDFFF0004020005D5555555A2AABFFFF5D516AA00A28028A00AAAEBF",
INIT_21 => X"3FEBA082ABFE10AAAEA8ABA55517FF45A2AEBDEBAAAAAA8BFFF7D140010FF841",
INIT_22 => X"FD75FF0051401FF5D00154105504000BA5D2E97545A28028B450855401450804",
INIT_23 => X"FBFFF45A2FFFDE00002E801FFA2AABFE00FFFFD74AA085540000002E801FF557",
INIT_24 => X"0000000000002ABEFAA80001EFF7FFC20BAF7D1575450800020BA08517FF45F7",
INIT_25 => X"57803AEBAF7F5D74AAA2A03AA38BF8FC00000000000000000000000000000000",
INIT_26 => X"7A3F00516DA2D5451D7EBDB47155BC2A87092AAFA9257F1C5BC00AA5D7FF8EAA",
INIT_27 => X"00EA8000150A801C01C7142EBFBC7EB8005B55A85B555EF095F50578085BE8FC",
INIT_28 => X"BEAE3D542A004380124921D20975FFAAA1521FF492BF8F40B6AAB84AF555168A",
INIT_29 => X"8F6DE05B40480557A95A3A1C2EBAE28168ABAA2D43D568BC5400168E90E2F412",
INIT_2A => X"47B50A80095178157FEFA0742FA3AA28EA8168A954100071D2E90A855C7A00A3",
INIT_2B => X"0A8F57F6DA971F8F7FFFA42D16D1EAE925EA0BFEBF4AA09217F4905684170851",
INIT_2C => X"000000000000000000000000000002D57AAA8402A8743DBD202DA95568A95E80",
INIT_2D => X"17D34ABA5D7BEAAAAD786BCEAAFFD1564BA2282BFA02A2C28000000000000000",
INIT_2E => X"007F8B2B2D97D483AFA7BD9F5EFA87F57555AAFBD7555FFAE95408A8FDC31AD0",
INIT_2F => X"0A6AEA8FAF0451CA001D4845C2087383F79A5046A37B55F38415555797D63BFF",
INIT_30 => X"A7D7463CC508D07577BAFBD542000D382964A92B401E71D7581C33172EC0A030",
INIT_31 => X"0502828811FCD4EABDB1DFDFC8365A2FD5E04AA5780A8AAAD7AC3CA02003BEBB",
INIT_32 => X"4FF72AAADF245595157050790621F562B1122DA70C3808458881056A5502AA15",
INIT_33 => X"F6A03D4BFB79AFA4C5CB5F5896D55BBAAC55EAFAF86D35E4A92B4460D1506037",
INIT_34 => X"FC0000007FC0000007FC0000007FC0000007FC0000007FC07AAF12E00505D3FD",
INIT_35 => X"7FC0000007FC0000007FC0000007FC0000007FC0000007FC0000007FC0000007",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000400000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"650C00000848A0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000004208B00200E010800006667BE7000102C00080000040012010000080C",
INIT_05 => X"0080000000002020600100208D04414000800000000200004800080000800200",
INIT_06 => X"04022140220932C2038900000100000008082010000000800488000000020400",
INIT_07 => X"088C0060242183060CF118011281B00000220010400020002081A00082100001",
INIT_08 => X"40000400014812466427040098C000622AAAA43E3060C158AC97F0356BDBFBD0",
INIT_09 => X"00026C000559102400200281400469000008B0800000901080004004308B4340",
INIT_0A => X"045413002200000000400408200000201041000208000040020820034200005C",
INIT_0B => X"41E11C008089540000420100101088400000808404004000000020A000100414",
INIT_0C => X"18C191AC191A4191A4191AC191AC191A4191A00C8560C8D08400000609010100",
INIT_0D => X"0E08A20BC417C16004C0B8382210904018000080100100012200000064064019",
INIT_0E => X"0E0615C96000000010200000802100022008100408020401020040100142200E",
INIT_0F => X"C06100000021E300B000000781E00140018000000781E00140018000002430E3",
INIT_10 => X"68C381C00000024E0000000781E00140018000000781E0014001908400005E11",
INIT_11 => X"088400003C30F00C000000155800D00000003E21C0700000000F001180000004",
INIT_12 => X"4000260640900004A400081401A0000004041218503E40300600000048043180",
INIT_13 => X"00009A0001208C30800025200003D807E0000000007252016000904618400013",
INIT_14 => X"480160000F00C0E06100000012D2005100409520381C00000005920004C0C812",
INIT_15 => X"0004025000120850B8180625400400000010711200510004B414780400000055",
INIT_16 => X"1004010040002002080000000804000A0000000011A000100208C008611430A0",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"5800050008000000000000000001004010040100401004010040100401004010",
INIT_1A => X"1451451451564090C69606492492C09A8C205148D757DF8A94102E0001063A29",
INIT_1B => X"BADD6EB75BADD6EB75BADD555555555555555555555555555555555555555145",
INIT_1C => X"FFE0000174BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974",
INIT_1D => X"F5D2AAAB555555400000000000000000000000000000000000000000000303FF",
INIT_1E => X"EFA2D17DEBAF7D1574BAAAFBFDFFFA2FFD74000855555FFFFFFC01FF087BE8BF",
INIT_1F => X"145557BFDEAA5500154AAAAAEBFF455D04175FF5D7FEAAAA002ABDEAA5D2EBFF",
INIT_20 => X"20BAAAD540145F7D5574BAAA8415400005540155F7D16AB45002EA8ABA005540",
INIT_21 => X"975EFF7AEBFF550055555FF55003DE00A2FFFFFEFAAD57DE00082AAAA00082A8",
INIT_22 => X"16AABAAAAEBFE10AAFBD7545F7D5554AA5D2ABDEBA082A821455D2EA8B455D2A",
INIT_23 => X"FFEABEFA2FBEAB455D7BD55FFFF84155FFFFFFFFF55AAAABFFFF5D556AB45A2D",
INIT_24 => X"000000000000175FFF7D140010FF84174BA552EBDEBA0004020AA5D04155FFAA",
INIT_25 => X"4BFBC51FF1471E8BEF55242FF47015A800000000000000000000000000000000",
INIT_26 => X"0B6AEBAEAA5D2EBDFFFBED17FEAAF7D5524AAA2F0BAF7FABDFC7E10005F525D7",
INIT_27 => X"55142A8708202FBD257F1C7550492490E17EAAA2AAB8F4515043DFC75575C700",
INIT_28 => X"03D1420AD000B420820AAE2DB6FB6DF7DFD5038ABA140A2D00554517DEBDB6FB",
INIT_29 => X"25555F8FFDE38087FC51C7F7AABFF55BC5B555C74B8A38E38085BE8B47A3A005",
INIT_2A => X"BA4AF555168B68FEDF6AB52AAABD21EF1C2FEA5FDEBDB505FA4920AFE10082E9",
INIT_2B => X"17AEB8BFF155552B6F5E8BFF1EFBFDBFF5FF1C00BF5D25475C7B7FEAFF45BEAA",
INIT_2C => X"00000000000000000000000000000151EAE3D542A004380124921D20BFFFA0AA",
INIT_2D => X"3D795000087BC01458AFBC11FF55516ABEFDD003EFE5093DC000000000000000",
INIT_2E => X"550434D555C53E0CE2AAA8742BA5D2ABDFFFF7D57DEAAFFD5420B2A2D37DB07A",
INIT_2F => X"F0851575FFAAFBDD5542B2EDD608897FD610D01151C610592A974BAFBAC28B55",
INIT_30 => X"100F3D68FFFAABAC20EF04003FE102400144ABAAFFF7DE772FDD56588042F72E",
INIT_31 => X"4EA0006BFE007E2E8315DD02F6A81A239501755F504BDF557D79431FD006EABA",
INIT_32 => X"03158517BD745AEAEA8FAF0C55EAF57FF957CAAA7FABF7DFD0C6A7DFFFA07FC0",
INIT_33 => X"964A92B403EE18D5408A6F2AFADF6900FFFF68BEFDFFB4B1FE5551141E78A028",
INIT_34 => X"0000000000000000000000000000000000000000000000165BAFBD542000D382",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000400000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0812",
INIT_01 => X"2145A00A1079284D04A044A54E504368404000720885800802000006ECD10200",
INIT_02 => X"5C010800020408040C415854AA055254090541A111000A104A00000009083510",
INIT_03 => X"0C1000100C0000D40526480250149120031500A0218808002440804288890550",
INIT_04 => X"8840C28120051400582012021808040409C0B26850488419444010C10A024A49",
INIT_05 => X"488510910548012025C0C0000300086854B141042252142042A048D090006372",
INIT_06 => X"948037480159A403109848000428AA8282102040449090D520085224410AA420",
INIT_07 => X"01020402242000408468112010810C055200022025A83AA3008882004A001542",
INIT_08 => X"11491C154429220A2824640010A010020282843E0008124C0000211000008840",
INIT_09 => X"E280442C1411D020828A2B116824632885419240016001900AE01A2020066395",
INIT_0A => X"30105108880684145002021012D40D718241108815380200900160AE42CE2818",
INIT_0B => X"53419F10308D100054AA080092112C100B400880454058E80B94080C49318000",
INIT_0C => X"D0090D0090D2890D0890D2890D0890D2090D0048610486808403A384880B8981",
INIT_0D => X"8202043800000620500403080A919000B8AD0304144008111A00582043243050",
INIT_0E => X"9835300002AA40AA902408200010002021060C810241832241280C81A0984020",
INIT_0F => X"100000000080A0000140000002000140200A8000000200014020100290E469C6",
INIT_10 => X"00100000000003400A8000000200014020094000000200014020087000000000",
INIT_11 => X"014200000004000000000081400004C00000000020000000008C000010A00000",
INIT_12 => X"0510000000000006800001880004008400800000000020000000000048100000",
INIT_13 => X"0000D0260000000000003409280000000000000040025000030000000000001A",
INIT_14 => X"400002A0000000000000000042900000A100000000000000008012A200000000",
INIT_15 => X"000000004420300000000000000000000010C010000098000000000000000105",
INIT_16 => X"00802208036408C0820010004D36A222120090554000E40080000000088000A0",
INIT_17 => X"8802008020080200822088220882208802008020080200822088220882208802",
INIT_18 => X"8320883200812008120081208832088320883200812008120082208822088220",
INIT_19 => X"E88051029FC0FC0FC1F81F81F820883208832088320081200812008120883208",
INIT_1A => X"08208208208C13A4301040B2CB2CBAC838B6C0080271AE180616A851158E2863",
INIT_1B => X"944A25128944A25128944A082082082082082082082082082082082082082082",
INIT_1C => X"FFE381F928944A25128944A25128944A25128944A25128944A25128944A25128",
INIT_1D => X"A550002000AA800000000000000000000000000000000000000000000003C200",
INIT_1E => X"BAFFAE801FF087BE8BFF5D7BEAA1055042AA105555421EFFFD568AAA002EBFEB",
INIT_1F => X"FFFA2D57DE10557BE8ABAF7AAA8BEFAAAE975FFA2D5555450851574000851554",
INIT_20 => X"5555F7D568ABAF7D5574BA552EA8AAA5D2EBFFFFA2D1554BAF7D17FEBAAAFFFD",
INIT_21 => X"EAAAA552AAAAAAAAAABFF455D04175FFFFD5574AAAAAA974BA082EA8BEFAAD55",
INIT_22 => X"FEAA000055401555D7BFFE10085557410F7AA97410087BD55FF087FEAA10A2FF",
INIT_23 => X"0017400550402155A2803FE005D7FE8B45F7FBFDE00085540155F7D56AA00007",
INIT_24 => X"00000000000017400082AAAA00082A820BAAAD540145F7D557410AA8428A1055",
INIT_25 => X"4BD16FAAA002ABFEAA550E82000E28A800000000000000000000000000000000",
INIT_26 => X"FEAFBD2410005F57482E3AA801FF1471E8BEF5574AFA00010ABFA38555F401D7",
INIT_27 => X"AAF7D5524AAA2F1FAF7FABFBFF400417FEF082F7AAA8BEFE2AA955EFA2DB5757",
INIT_28 => X"492082EADBFFBEDB55555E3DF6DA82F7DF520385D2FE80AA5D2EBDFD7BED1574",
INIT_29 => X"21C7005B6FB47F7A438E925D24ADAAAB6AAB8F455784155C75575C7000B6AE95",
INIT_2A => X"4717DEBDB6FA3D0075EDA800051C05571474024A81C5557578EBA087400007FC",
INIT_2B => X"FFDE381D716FA15550015428E10A001FFB40038F68F7F578F7FFEF568E280855",
INIT_2C => X"000000000000000000000000000001043D1420AD000B420820AAE2DB4716DF7D",
INIT_2D => X"828FDEBA5D7BC015582D57DEAA002ABDEAA552A80010AAA88000000000000000",
INIT_2E => X"AAAE955EFAAFBC15F5A3D7D6800087BD5410AAAA801FF55556ABEF5D517EEE00",
INIT_2F => X"A5D2ABDF55F7D575EAAFFD50A2B2A3D169B07A3D7BFE10597BFDE00AEAC28BFF",
INIT_30 => X"555A53C00B2A2AA02000082ABDFEFFFFBC1154AAFFFFE107FF9D72A20842080B",
INIT_31 => X"4EAA28015400547FC315D00797CF4780286A2105D2A3FEBAFFAC28B555504145",
INIT_32 => X"99ADABD5A8AAA0051575FFA2FFFDA02003FFDEAA8557D65550915544AA5D5157",
INIT_33 => X"144ABAAFFD75E7F2BDDD2B8016F9E2555500174AA282E20BFFFF842AAAAADD56",
INIT_34 => X"0000000000000000000000000000000000000000000000030EF04003FE102400",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000800000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380206",
INIT_01 => X"200C9A40408001683C0462C99E004B61404040028804A0080A000416A0990A0C",
INIT_02 => X"4809A900031800444461089866E331352180D468B8040E600C0081110B802CD0",
INIT_03 => X"6D0B61108C00014231A3080408C68420330066010A80881068A808401CC46330",
INIT_04 => X"482218066A09C03B348C1C1928DD5A4402211A68470944842640902107002D24",
INIT_05 => X"0583180353202020000144E50B44644B30A86D05014A0D224063095092100E34",
INIT_06 => X"54023740216934020303680A040066D98A182210085A50C02048288234629414",
INIT_07 => X"018C00220430814204E01C581291820CCA000E3226413990008C80205A00CCCC",
INIT_08 => X"4108747320081246252D5010184000220002A43E10294258E805E1156002D940",
INIT_09 => X"D0AA546AC41B112029A61D84424429AA1320B1010140C1350B48292020024180",
INIT_0A => X"000102022850A1CC0047071913208CE802430488082042008040F399606F4058",
INIT_0B => X"5141BE42B88840005268081412152900484201A814144D60888CAA2C48151020",
INIT_0C => X"1B49019490194901B4901B4901949019C901B64805E480CA94480506980125C4",
INIT_0D => X"5A01E2B1080602E00C54216800859000199C98800C8140A11A44423040240450",
INIT_0E => X"28A65300E6664599902600009821204A040C1C040C0205038300480801480208",
INIT_0F => X"000000000090000003202900000010002008A02900000010002008039666928B",
INIT_10 => X"00000000000801000A202900000010002009E0290000001000200A3800008000",
INIT_11 => X"036000008000000000000088000002D003008000000000000280100016200812",
INIT_12 => X"05B008088000008201021C880000488002810005000000000000040000100000",
INIT_13 => X"0010402B80412000000410199800040000000000408020000680209000000208",
INIT_14 => X"800012980040300000000000C020000C8300208800000000008200AE01011000",
INIT_15 => X"40A0000841003100010401000000000002008020000C38000200000000000120",
INIT_16 => X"10070300704028820801400068360424820185CCE0128010020000008088021C",
INIT_17 => X"0070100701007010050180501805018050180501805018070100701007010070",
INIT_18 => X"070140601007014060100701C040180501C040180501C0401807010070100701",
INIT_19 => X"4A81454A26AA555AAB554AAB5541C040180501C040180501C040180501406010",
INIT_1A => X"08208208209441D0B0000092492480AA2860607818F18E0C851428200B262C31",
INIT_1B => X"D4EA753A9D4EA753A9D4EA492492492492492492492492492492492492492082",
INIT_1C => X"FFD55E21A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8",
INIT_1D => X"FAA8000155080000000000000000000000000000000000000000000000000200",
INIT_1E => X"EFFFD568AAA002EBFEBA555142000AA802AA10F7D57FEAA557BE8B45A2D5555E",
INIT_1F => X"A10550402000AAD56AAAA557BC0155A280021EFA2FFE8B4555042AA105555421",
INIT_20 => X"0010AA842AAAAFFD542000FFD5574000851554AAFFAE801FF087BC01FF5D7FEA",
INIT_21 => X"7DE105551420BAF7AAA8BEFAAAE975FF005540145A2D157410AAD17DFFF5D040",
INIT_22 => X"03DEBAAAFFFDFEFAAD57DEAAF7AE975FF080428B455D7FFDEAA5D55574BA0051",
INIT_23 => X"AE800AA087BD5555552A821EF007FFFEAAAAD5554AA552EBFFFFA2D5554BAF78",
INIT_24 => X"000000000000020BA082EA8BEFAAD555555F7D568ABAF7D5574BA552E800BAAA",
INIT_25 => X"E975EAB6DBEDF575FFAA8E02155080E800000000000000000000000000000000",
INIT_26 => X"5EBAEADA38555F451D7EBD16FAAA002ABFEAA555E02000E28AA8A38EBD578E82",
INIT_27 => X"FF1471E8BEF5575EFA00012A87A38AAD56DA824975C217DAA84021FFAAF5EAB5",
INIT_28 => X"400BED57FFD7410E05038BE8E2DABAFFDB47412ABFE90410005F57482E3AA801",
INIT_29 => X"FEBA5D71D742A407FFFE00555F47082E3AAA8BEFA02A955EFA2DB5757FEAFBD2",
INIT_2A => X"BFFD7BED157482F7803AEAAA2F1FAF7FABFBEAE2AEBA4974871C043AB6D4975F",
INIT_2B => X"F7AE38497FC00BAB6A4850821C75D25C74920821D708757AE2AA3FFC04AA552E",
INIT_2C => X"0000000000000000000000000000007092082EADBFFBEDB55555E3DF6DA82F7D",
INIT_2D => X"AA8A8ABAAAD568A1020516ABFFFFFFD75FFAAAE8014500288000000000000000",
INIT_2E => X"AA80001FFAAD57EB55A2A8ABEBA5D7BD5545A2D57DEAA002EBDEAA557BC0010A",
INIT_2F => X"0087BD5410AAAA801FF5555629EF5C517EEE00828D74AAFBD57DE000057C21FF",
INIT_30 => X"EFA8FBC15E5A3D5D7400FFD57DF55082E974AAFFAABDEBA77FDD66A0ABBDC200",
INIT_31 => X"50555002ABFF54517EEB25D57C14100957FF6105D7BD5400AAAC28BFFAAAE955",
INIT_32 => X"FA42A3D7020BA5D2ABDF55F7D1554A8FFC42AA10A7D169F57ABD7FEEBAAA8415",
INIT_33 => X"C1154AAFFFFE10FFF9DF202096F014AAFF84154105555C215500000014558557",
INIT_34 => X"000000000000000000000000000000000000000000000015400082ABDFEFFFFB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000400000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204002",
INIT_01 => X"01039802000820491C00650E1E004340403008418984014902030906A8D10200",
INIT_02 => X"480108A000000000444048E41E80F00A41043118680002000800000009882390",
INIT_03 => X"06504110080000D0040608024010102026001260300000003080880208C000F0",
INIT_04 => X"9100E98268154C1AE0B01C160033B944028290285AE0DC38E02090E81C22E801",
INIT_05 => X"5C0F20B36F000109200044C401041C4CF21C48B433483C8242EAE1B0000074C4",
INIT_06 => X"100007000059800310086A1A0022E18780000140C9D9D0930000F228075A6071",
INIT_07 => X"00000000242000008461000810818403C100060064012E00048C82201800BC28",
INIT_08 => X"0048CC8F01090602202C0400008000002202243E400010480000211540008810",
INIT_09 => X"40E0DC1EB5191120C7BE7D152201612E80E891E0614041340838450020422111",
INIT_0A => X"30545DAD8C2E0982400603003200872003FB1408082840002044007846164E0A",
INIT_0B => X"43411D10118D1A04522E000498140C104B260DA0404003C08B6000AC01128000",
INIT_0C => X"C5010C3010C1010C3010C1010C1010C3010C140869808618850BE6305989AB80",
INIT_0D => X"100140302800108018840440028480001B8780800000003102045C3443043410",
INIT_0E => X"3080620481E0E18790012A001001026808000002020101028100200180080201",
INIT_0F => X"000000000010000005C0200000001000000C4020000000100000000380E4C308",
INIT_10 => X"00000000000800000D00200000001000000EC020000000100000086A20008000",
INIT_11 => X"012820008000000000000008000001B00100000000000000020000002AA00010",
INIT_12 => X"06D0000080000080000241D80000800442800001000000000000040000000000",
INIT_13 => X"0010003A00002000000400021800040000000000008010000B00001000000200",
INIT_14 => X"400005900000100000000000801000089000008000000000000200F800001000",
INIT_15 => X"00000000A500100000000100000000000200001000002E000200000000000020",
INIT_16 => X"000000C032700000022400444934240A8021B63C005108010004100098098010",
INIT_17 => X"C010080200401008000040300800004010000200C01000020040100802004030",
INIT_18 => X"02000000000100C0300400008000000300C0100C00000020080000C030000000",
INIT_19 => X"20240142325930C9A6CB261934C000200801004030040200800000030040100C",
INIT_1A => X"14514514514E98264686668A28A260521CC45140C700FC0A0002870980831A28",
INIT_1B => X"1A8D46A351A8D46A351A8D555555555555555555555555555555555555555145",
INIT_1C => X"FFD5E7D8341A0D068341A0D068341A0D068341A0D068341A0D068341A0D06834",
INIT_1D => X"A5D55420AA002A80000000000000000000000000000000000000000000000200",
INIT_1E => X"AA557BE8B45A2D5555EFAAD140155080000155FF843FFEFAA84001FF5D043FEA",
INIT_1F => X"000AA80001555D04174AA002A80010FFAE975FFAA80001EFA2AAAAA10F7D57FE",
INIT_20 => X"00BA5D51555EF002AA8BFFAAAAAAA105555421EFFFD568AAA002EBFEBA555542",
INIT_21 => X"82000AAD568AAA557BC0155A280021EFA2FFE8B45F78400145FF842AAAAA2AA8",
INIT_22 => X"BC01FF5D7FEAA105D0428B4500003DFEF080428B455D002AABA5D2AAAAAA5D2E",
INIT_23 => X"80154BAA2FBE8AAAF7AA821EFAAAAA8BEF552E820000851554AAFFAA801FF087",
INIT_24 => X"00000000000015410AAD17DFFF5D0400010AA842AAAAFFD542000FFD57DF55A2",
INIT_25 => X"A284051D755003DE92415F42092142E000000000000000000000000000000000",
INIT_26 => X"71C0A28A38EBD57DE824975EAB6DBEDF575FFAADE02155080E85145E3803FFEF",
INIT_27 => X"AA002ABFEAA555F42000E2AA851455D0A124BA002080010FFA4955C7BE8E021C",
INIT_28 => X"145F7802AABAA2A480092415B505D71424AABD7F68E2FA38555F451D7EBD16FA",
INIT_29 => X"AA824924AAA92550A07038BED56DA824975C217DAA84021FFAAF5EAB55EBAE82",
INIT_2A => X"55482E3AA801FF1471C01EF5575EFA00012ABFB6D080A3AFEF080A2FB45490E2",
INIT_2B => X"B6FA12ABAEBDF7DAA80104BAAAFFEAA00F7AE821D7B6A02FBC71D0E10010005F",
INIT_2C => X"0000000000000000000000000000010400BED57FFD7410E05038BE8E2DABAFFD",
INIT_2D => X"02897555A2803FFFFAA841754555043FE10087BC2000552C8000000000000000",
INIT_2E => X"FF8017545F7AE821455D2CAAABAAAD57DE1000516ABFFFFFBD75FFAAFFC01450",
INIT_2F => X"A5D7BD5545A2D57DEAA002EBDEAA557BC0010AAA895555042E820BA080400010",
INIT_30 => X"FFAAD57EB55A2A880155F7802AAAAAA8002010007FC0155D5022A955FFACBFEB",
INIT_31 => X"BEF002EBDF45542AAAA0008043CAB0552C97CAAFFD57DE000057C21FFAA80001",
INIT_32 => X"CFE55D2CC2000087BD5410AAAA801FF5555421EF58517EAB00028A9BEF002EAA",
INIT_33 => X"974AAFFAABDEBAF7FDDE6A0AA90FDFEFA280020BAA2FFEAA10FFAE82145F7803",
INIT_34 => X"000000000000000000000000000000000000000000000002000FFD57DF55082E",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000800000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A337A20E07C0C1E006",
INIT_01 => X"295FBC468000A04D5C6A60000C34C24841280A00084000C8C212892EEAD53235",
INIT_02 => X"C809AD5CB118E640A4D158F8011FF0002080000082C8C66609DB7DDDCB1F2036",
INIT_03 => X"250906263A4C904214A35C80085285720B20648A88800000B8E0F852A884500E",
INIT_04 => X"4005122126899100064D20001044429C78A43A2C4436CC87198A3916E0551A24",
INIT_05 => X"A370C14CA0E900004048402389CFE2F20F7D7A354CB5C208E51437F044948912",
INIT_06 => X"9B9407B9424F33468B096FCF452AE0505A185905CC2414D44437118630839B88",
INIT_07 => X"588C732074A68D5AB4EB180717FF513FC52691924098712CE481FDC201D43C1A",
INIT_08 => X"0016053F180A1286A4ED1BC18840C320000055FE91AA545CBA4DE1D17992D9BE",
INIT_09 => X"2D1A4D8105B734723041008100486100601EDE1DE46431138DFD404CB4022595",
INIT_0A => X"A131112C0D15C901B2122309204C28B67061E81A8920C8D3CF8014007902DA6B",
INIT_0B => X"AD5C3402488888E5126BA350B27C092E63D18C9C500577EEA33EF24C09B42464",
INIT_0C => X"096B80D6B80B6B80F6B8096B80F6B80B6B80D15C04B5C07AD50C94020D233107",
INIT_0D => X"8948020D829FA454104132252011E542387F810480C840C383751EF5606E0178",
INIT_0E => X"000200CA7FE0627FD25845E42151648F854480A042512028100A8C38280AA04C",
INIT_0F => X"D06101C55DE5E3E3C017E37FC3E0017C3F8817E37FC3E0017C3F900040241001",
INIT_10 => X"6CD381C0118797FE0817EA7FC3E0017C3F8817EA7FC3E0017C3F9900DFFFDE15",
INIT_11 => X"F800DFFFBE34F00C0270F3F55F1F8007FDBEBE25E0700463E1FF2C7E014FF7BE",
INIT_12 => X"C5DEF64EC090626FE40140459759173BBD6EF37D523E6030061341F07FD571F8",
INIT_13 => X"0C4DFE2A6FE2AC3082637F281BFFFC07E00007E07F7253D38337D1D6184131BF",
INIT_14 => X"4F4F8397FFA0F0E06101C53E76D3D3E884FDDDA8381C0098E5FD92BBDFC8D812",
INIT_15 => X"19074FA36FDF58DBF81C072540049707E0FEF313D3E03BFFF61478040570EFD5",
INIT_16 => X"8CA02ACA00C50850182309444D248204201040FC190054A2110B8ACC483204A1",
INIT_17 => X"0A128CA0284A2280A1288A128CA2284A0288A1288A3284A228CA0288A1280A32",
INIT_18 => X"A228CA0284A3280A3288A1288A3280A2284A028CA2284A2284A028CA0280A328",
INIT_19 => X"F6A1850E1892596D34924B2DA6A84A2284A1288A1280A3280A1288A0284A2284",
INIT_1A => X"7DF7DF7DF7CBFBFE7EFEEE79E79EFAF3F51EB769CFEF73B6FFE74FC2400DB6DB",
INIT_1B => X"EEF77BBDDEEF77BBDDEEF77DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF",
INIT_1C => X"FFC27F6BDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDD",
INIT_1D => X"55D2E955FFF7FFC0000000000000000000000000000000000000000000000200",
INIT_1E => X"EFAA84001FF5D043FEAA5D04020AA002AAAABA555140155087FFFFEF00042AB5",
INIT_1F => X"1550800001FF5D00001555D2E975FF5D5568B555D7BD5545FFD540155FF843FF",
INIT_20 => X"FF45A2FFC0000AAAE974AAFFFFEAA10F7D57FEAA557BE8B45A2D5555EFAAD540",
INIT_21 => X"401555D04174AA002A80010FFAE975FFAA80001EF002AAAABAF7D168A10A2D17",
INIT_22 => X"EBFEBA555542000A28028BFFF7803DF55FFAEBFE005D2EAAB45557BD55555555",
INIT_23 => X"517DF55082E974BA087FE8B55552E955EF5D7FEAA105555421EFFFD568AAA002",
INIT_24 => X"00000000000000145FF842AAAAA2AA800BA5D51555EF002AA8BFFAAAA820AA5D",
INIT_25 => X"007FFFFFF1C042FB7D492A955C7F7FBC00000000000000000000000000000000",
INIT_26 => X"5E3DB45145E3803AFEFA284051D755003DE92410F42092142E28ABA5D5B4516D",
INIT_27 => X"6DBEDF575FFAADF42155082E851C75D0E02145492E955C75D5F6DB55497BD554",
INIT_28 => X"ABAF7D16DA28A2DB7AF7DB6FBC7028A2AA95492FFFFE8A38EBD57DE824975EAB",
INIT_29 => X"FB45557BD5555415F45145490A124BA002080010FFA4955C7BE8E021C71C0A2D",
INIT_2A => X"451D7EBD16FAAA002ABFEAA555F42000E2AAA8BEFE3843AF55E3AABFE105520A",
INIT_2B => X"4821D7F68E07082495B7FF7D082E954AA087FEDB7D5D2A155D7157BEFA38555F",
INIT_2C => X"0000000000000000000000000000002145F7802AABAA2A480092415B505D7142",
INIT_2D => X"52CAAAAA5D7FD75EF087BFDFEF5D003DFEF002E95555F7FDC000000000000000",
INIT_2E => X"5D7BFDF45007FD7555A2F9D5555A2802ABFFAA841754555043FE10082A820005",
INIT_2F => X"AAAD57DE1000516ABFFFFFBD75FFAAFFC0145002895545552E80145002E95545",
INIT_30 => X"45F7AE821455D2CBFEAAFFD17FEAAAAFFEABFFF7FFD54BAA2AA95410F7FDEAAB",
INIT_31 => X"B45AAAABFE0009043FF555D7BD55550879D5555002E820BA080400010FF80175",
INIT_32 => X"75455D7DFFEBA5D7BD5545A2D57DEAA002EBDEAA557BC0000AAA8A8BEFA28028",
INIT_33 => X"02010007FC0155550222955FFAC97400087FFFFFF002E954AA087BFFFFF5D2E9",
INIT_34 => X"000000000000000000000000000000000000000000000000155F7802AAAAAA80",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000003000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B0061A258A2840112C03002C180004003220200403302301C0381A0086",
INIT_01 => X"860041C83839484C00A100000052024841000000090800090210010000510204",
INIT_02 => X"080108200C1000004464080400C0080100000000010432400800800009882050",
INIT_03 => X"040001008C2340D0800208624200002183800584488000103080010C08C10000",
INIT_04 => X"00101610A029B08400044800000000040008102A040810040400900500001800",
INIT_05 => X"02800000400C830934E4A0002900404400820000000A00824004084011200A00",
INIT_06 => X"14C8874C884D0C024608680210C11F8010122100880802800308010000829400",
INIT_07 => X"060800002430200004611000508184803A0900224000200008818028C04883E1",
INIT_08 => X"4041FE80E009024260240010608000000000043E040000488000201400008810",
INIT_09 => X"0002447E041B112020208010404029006FE0B081003204502000002068621191",
INIT_0A => X"35E5148B0D916BBE39049191200000200441048108000220002FC5FA60000148",
INIT_0B => X"5358BF12E88D1000022808801A112D1443142A815440600083FE9AA300100281",
INIT_0C => X"C1416C1416C5416C5416C3416C3416C7416C500B60A0B60AD40E34104C093904",
INIT_0D => X"8C03403C440C054048850A300A8480009A0020865AE4ECB11B441A105B05B016",
INIT_0E => X"00000031001E4800022100321489214001A742D3A368D1B4686D100234B44242",
INIT_0F => X"00000000000AB800302008000000014000602008000000014000674000260000",
INIT_10 => X"0000000000000241E020010000000140006020010000000140006A8400000000",
INIT_11 => X"028400000000000000000003C00052000200000000000000000CD00184000800",
INIT_12 => X"30000800000000049A48184000A0400000010000000000000000000048028C00",
INIT_13 => X"0000918480010000000024C9E000000000000000000FF0006440200000000012",
INIT_14 => X"C000602800400000000000000BB000112B0020000000000000007E0000010000",
INIT_15 => X"02A0005000202500010000000000000000104CF000198000000000000000000F",
INIT_16 => X"4AD2B46D180684E8402440044C24A30819020603E0A20640C8400010218432A0",
INIT_17 => X"2D1B4ED3B4AD0B42D1B4ED2B42D0B46D1B4ED2B42D1B46D3B4AD2B42D1B46D2B",
INIT_18 => X"D1B42D0B46D2B4AD1B46D0B4AD3B4ED0B46D1B4AD2B4ED1B42D0B4ED3B4ED0B4",
INIT_19 => X"F8840000331C618E38E38C31C7346D3B4AD3B46D0B42D3B4ED2B42D1B42D2B4E",
INIT_1A => X"1C71C71C71CEDBB676F66EFBEFBEFAF99CFEF179CFF1FE1E9F52AFF9BFAFBE7B",
INIT_1B => X"FE7F3F9FCFE7F3F9FCFE7F1C71C71C71C71C71C71C71C71C71C71C71C71C71C7",
INIT_1C => X"FFE43591FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"05D2EBDF55557FC0000000000000000000000000000000000000000000030200",
INIT_1E => X"55087FFFFEF00042AB555D2E955FFF7FFC21EFF7D17DEAA5D2AAAAAA5D557DE1",
INIT_1F => X"0AA002A82145555542010FF803DEAA5D5568BEF5D042AA10A2AAAAABA5551401",
INIT_20 => X"20BA00557DF455D7BFFEAA555540155FF843FFEFAA84001FF5D043FEAA5D0002",
INIT_21 => X"001FF5D00001555D2E975FF5D5568B555D7BD5545FFD568AAA5D00154AAAAD14",
INIT_22 => X"5555EFAAD540155080000000F7843FF55007FFDEAAA284020BAAAD168BFF0800",
INIT_23 => X"51401EFF7842AA00FF8417545AAAEBFE10FFFFEAA10F7D57FEAA557BE8B45A2D",
INIT_24 => X"0000000000002AABAF7D168A10A2D17FF45A2FFC0000AAAE974AAFFFFC21EF55",
INIT_25 => X"5520ADA92495B7AE10412EBFF45497FC00000000000000000000000000000000",
INIT_26 => X"0AAAAA8ABA5D5B4516D007FFFFFF1C042FB7D492A955C7F7FBC71EFFFD57FE82",
INIT_27 => X"D755003DE92410E02092140E0716D415F47000F78A3DE92415F6ABD7490A28A1",
INIT_28 => X"A92550A104AABED1470AA005F78F7D497FFFE925D5B45145E3803AFEFA284051",
INIT_29 => X"20BAA2DB68BC7140E051C75D0E02145492E955C75D5F6DB55497BD5545E3DB6A",
INIT_2A => X"7DE824975EAB6DBEDF575FFAADF42155082E87038FF8038F6D1C7BF8EAAAA800",
INIT_2B => X"A95492FFFFC71EF415F471C7FF8428A00E38412545AAAE3FE10A3FBE8A38EBD5",
INIT_2C => X"000000000000000000000000000002DABAF7D16DA28A2DB7AF7DB6FBC7028A2A",
INIT_2D => X"7FDD55EFF7D57DE005D003DE00007FEAA10002ABFF450079C000000000000000",
INIT_2E => X"087BE8B45082EAAA10A2A8AAAAA5D7FD75EF087BFDFEF5D003DFEF002E95555F",
INIT_2F => X"5A2802ABFFAA841754555043FE10082A82000552C955FF007BD5410FFAABFE00",
INIT_30 => X"45007FD7555A2F9EAA005D2A820AAF7D5574AA087BEABEF007FFDE00557DD555",
INIT_31 => X"BFF557BE8ABAA284020BAA2FBEAB55552C95545552E80145002E955455D7BFDF",
INIT_32 => X"FE10A2F9EAABAAAD57DE1000516ABFFFFFBD75FFAAFFC01450028974BAFF842A",
INIT_33 => X"EABFFF7FFD54BAA2AA95410F7FDD55EF007BD5555F7802AA10AA8000145AAAEB",
INIT_34 => X"00000000000000000000000000000000000000000000003FEAAFFD17FEAAAAFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000002400000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0048201002842002C02450018800002300500030B313300C418992002",
INIT_01 => X"A34009C23838684D1C20E0000E11426840000000080000080200080000110200",
INIT_02 => X"4801082048100000446558040080000041000000000622400800000009000010",
INIT_03 => X"040001818CA144D0842248424210812103000480088000003080014688800000",
INIT_04 => X"000012002041900000048000000000040088322944200C850001940400301800",
INIT_05 => X"0200000040084000284000204104004402000025000800065004207030320800",
INIT_06 => X"108017080149000246086A2A1468004012120004440812D40120008200829001",
INIT_07 => X"2408000024302040846810005281848003494020400031240C8C8218E06A0009",
INIT_08 => X"4040050001090242602C0418408000000000243E0408104C8000201540008810",
INIT_09 => X"00024401041B132820000001424069004000B204636009104A0101226A422104",
INIT_0A => X"80049800A0281400300B0210200008B206639389480046240068180262000048",
INIT_0B => X"41401C1081811C44D22A18841616004118004482040448011800004D49340082",
INIT_0C => X"00192001920019200192041920419204192060C9010C90100008040008012101",
INIT_0D => X"48A000880144434A001001228000803198003604004048294008C40C483480D2",
INIT_0E => X"0000002160006000100000200811020805000480004000220108000060000800",
INIT_0F => X"09864038A2881210382000000001E003E0582000000001E003E0422834240000",
INIT_10 => X"0000160700706901982000000001E003E0582000000001E003E04E8400000000",
INIT_11 => X"0684000000000330C00F0C8210807200000000000581C01C1C809201C4000000",
INIT_12 => X"29D000000C2419121028C00020A2400000000000080082C180603A0E003A0904",
INIT_13 => X"8322414E800000432118908DF8000000061E001FC00C10207740000021908C48",
INIT_14 => X"40806BB800000009864038C14810201BAB000000026130071A80613A00000184",
INIT_15 => X"840080546520350000600812058100F81C018890201BBA0000008239020F1108",
INIT_16 => X"04812208033400C0022140404D268624B210040004A08400000044222900320C",
INIT_17 => X"0832048120481204822008020080204832048120480200802008020081204812",
INIT_18 => X"802008020C812048020080200812048120080200802048120483200802008020",
INIT_19 => X"0221054A2C208200010410400020880200812048120C80200802008120C81200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFD3B3D800000000000000000000000000000000000000000000000000000000",
INIT_1D => X"5AA8017410555540000000000000000000000000000000000000000000000200",
INIT_1E => X"AA5D2AAAAAA5D557DE105D2EBDF55557FFDE00557BEAABAA2AEAABEFF7801555",
INIT_1F => X"5FFF7FFD5555557BEABFFF7FBEAAAAAAD157555AA803FEBA5555421EFF7D17DE",
INIT_20 => X"DFEFAA80000BAAAAA820BAA2802AABA555140155087FFFFEF00042AB555D2E95",
INIT_21 => X"02145555542010FF803DEAA5D5568BEF5D042AA10A2AA955EFF7FFD5400F7FFF",
INIT_22 => X"43FEAA5D00020AA002ABDEBA5D7FE8A000004154BAF780001EFAAAAA8B450000",
INIT_23 => X"2AAABFF5551421FFAAD157545AAD5555EF557FC0155FF843FFEFAA84001FF5D0",
INIT_24 => X"00000000000028AAA5D00154AAAAD1420BA00557DF455D7BFFEAA5555575455D",
INIT_25 => X"AAA0A8BC7EB8417555AA84104385D55400000000000000000000000000000000",
INIT_26 => X"A4155471EFFFD57FE825520ADA92495B7AE10412EBFF45497FFFE385D71E8AAA",
INIT_27 => X"FF1C042FB7D492A955C7F7FBD056D5D75EABC7FFF5EAAAABEDF5257DAA8438EB",
INIT_28 => X"5EFEBFFD2400EBFBFAFEFAA80070BAA2A0870BAAA8028ABA5D5B4516D007FFFF",
INIT_29 => X"01D7AAA0AFB6D1C040716D415F47000F78A3DE92415F6ABD7490A28A10AAAA92",
INIT_2A => X"3AFEFA284051D755003DE92410E02092140E3DE924171E8A281C0E10482F7840",
INIT_2B => X"FFFE925D5B525454124AFBC74955421EFA2DF5557DAAD5D05EF0175C5145E380",
INIT_2C => X"000000000000000000000000000002AA92550A104AABED1470AA005F78F7D497",
INIT_2D => X"079FFEAA5D5568ABAA2842AB55A28015545A284000BA5D534000000000000000",
INIT_2E => X"F7FBC01EFA2842AABA0857555EFF7D57DE005D003DE00007FEAA10002ABFF450",
INIT_2F => X"A5D7FD75EF087BFDFEF5D003DFEF002E95555F7FDC01EF55556AB55F7D56AABA",
INIT_30 => X"45082EAAA10A2A8801FFA2FFC2000A2FFEABFFAA84174BAAA80174AAAA862AAA",
INIT_31 => X"AAA552A80010F78000145AA843DFEF5D02155FF007BD5410FFAABFE00087BE8B",
INIT_32 => X"21FF085755555A2802ABFFAA841754555043FE10082A82000552CBFE10085168",
INIT_33 => X"574AA087BEABEF007FFDE00557DC014500003FF450051401FFA2FBD55EFAAD54",
INIT_34 => X"00000000000000000000000000000000000000000000002AA005D2A820AAF7D5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"A14008420008204D042100000212026840000000180800080200090048510204",
INIT_02 => X"080108000090000004655C040080000051000000000402400800000009000010",
INIT_03 => X"00000100803008D0842240024210810003800584488000103080894288800000",
INIT_04 => X"00009610A028B084000440C0040000040088323244280C950400808500321800",
INIT_05 => X"42800080400C8A09306420202804400402800035200A00020204287001114A00",
INIT_06 => X"14C8864C8849880002486800142BFF001292214444081254002801A200821400",
INIT_07 => X"004800002430204084281000D281040001182020400031241C0D80000041BFE9",
INIT_08 => X"444005000108020220240010048000000000043E0408104C8000000100008810",
INIT_09 => X"0812040105191100200081130210ED104008A285617205D02A01010141225091",
INIT_0A => X"8004C8252291490039039390200008B20E230008280040088040100240008061",
INIT_0B => X"40013C128BC95C44522A00241204094008442681100448000800826F49240001",
INIT_0C => X"0408000080000800008000080000800008000440020400229548040008012125",
INIT_0D => X"401140BC4028430108150900408590109A00209642E46CA00240460400200440",
INIT_0E => X"080410010000200002210A320C89000005A142D0A16850B6294D100234201242",
INIT_0F => X"2F9EC00000800008100020003C1FE00020080020003C1FE00020044014260082",
INIT_10 => X"132C7E3F00000100080020003C1FE00020080020003C1FE000200880000081EA",
INIT_11 => X"0080000081CB0FF3C000008000201000010001DA1F8FC0000080110080000010",
INIT_12 => X"040000B0BE6C00020040580040200000001004832CC19FCF81E0000000100002",
INIT_13 => X"80004020000C31CF60001000000007F01FFE00004000300420000618E7B00008",
INIT_14 => X"C0102000000F151F9EC0000040300401000200D547E3F00000800080001617AD",
INIT_15 => X"02A020100000822406E1B95A3F83000000008030040100000BAB87FB00000100",
INIT_16 => X"46D1B66D1A368C68D26000544D26A504AB120400222206404840001101843000",
INIT_17 => X"2D1B46D1B46D1B46D1B46D1B46D1B42D0B42D0B42D0B42D0B42D0B42D1B46D1B",
INIT_18 => X"D1B46D1B42D0B42D0B42D0B42D1B46D1B46D1B46D1B42D0B42D0B42D0B42D0B4",
INIT_19 => X"20840442200000000000000000346D1B46D0B42D0B42D0B42D0B42D1B46D1B46",
INIT_1A => X"3CF3CF3CF3DBF91E66C6FAD96D965201F4C251414A87D78AF421448BE28F3AEB",
INIT_1B => X"3E1F0F87C3E1F0F87C3E1F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"FFD160B27C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C",
INIT_1D => X"AFFFFC2000557FC0000000000000000000000000000000000000000000000200",
INIT_1E => X"BAA2AEAABEFF78015555AA80174105555420000000021EFAA843DE00F7803FEB",
INIT_1F => X"F55557FD54AAA2AA955FF00043DE005504175FF08514014555557DE00557BEAA",
INIT_20 => X"DF45FFD17DFFFFFD56AA00557FC21EFF7D17DEAA5D2AAAAAA5D557DE105D2EBD",
INIT_21 => X"55555557BEABFFF7FBEAAAAAAD157555AA803FEBA55556ABFFA280154BAFF803",
INIT_22 => X"42AB555D2E955FFF7FFD5410002AAAAAAA2D57DF450004154BA087BEAAAAF7D5",
INIT_23 => X"843DE1008556AA00A28028B55FFD1555EFA2802AABA555140155087FFFFEF000",
INIT_24 => X"000000000000155EFF7FFD5400F7FFFDFEFAA80000BAAAAA820BAA280000AAA2",
INIT_25 => X"A2803AE38FF843DEBAEBFFC20285D75C00000000000000000000000000000000",
INIT_26 => X"55D5F7FE385D71E8AAAAAA0A8BC7EB8417555AA84104385D5542038000A001C7",
INIT_27 => X"92495B7AE10412EBFF45497FD24BAA2AA955C708003FE285D00155FF00554515",
INIT_28 => X"BEFA28E124AAF7843AF7DEBDB78FFFE3DF6DA284175C71EFFFD57FE825520ADA",
INIT_29 => X"04920875EAA82F7DB5056D5D75EABC7FFF5EAAAABEDF5257DAA8438EBA415568",
INIT_2A => X"4516D007FFFFFF1C042FB7D492A955C7F7FBD54380020ADA82BED57DF4508041",
INIT_2B => X"0870BAAA80070BAA2803DE00005F68A10BE802DB55E3DB555FFF68028ABA5D5B",
INIT_2C => X"00000000000000000000000000000125EFEBFFD2400EBFBFAFEFAA80070BAA2A",
INIT_2D => X"D53420BA082E82155AA802AAAAFF803DEBAAAFBC20BA55514000000000000000",
INIT_2E => X"5D04175EF0855575455D7BFFEAA5D5568ABAA2842AB55A28015545A284000BA5",
INIT_2F => X"FF7D57DE005D003DE00007FEAA10002ABFF450079C20BAAAAE9754500043DEBA",
INIT_30 => X"EFA2842AABA085768BFFA2AE820AAFF802ABEFAAFFEABEFAAFFFDEAA0051555E",
INIT_31 => X"E10F7D17FF5500000001008516AA10FFFFC01EF55556AB55F7D56AABAF7FBC01",
INIT_32 => X"75EFF7842AAAA5D7FD75EF087BFDFEF5D003DFEF002E95555F7FDD74BA08043D",
INIT_33 => X"EABFFAA84174BAAA80174AAAA86174AAAA843DE00087FE8A00F7843FF45AAFFD",
INIT_34 => X"0000000000000000000000000000000000000000000000001FFA2FFC2000A2FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000001000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"A1400802000020490000000000000240413C0A61590001D90213C90008510204",
INIT_02 => X"680108200010000054655C040080000041000000010402400800800009082011",
INIT_03 => X"00040100800020D0842240124210810043800504488000103081894288800000",
INIT_04 => X"00001410A00AA084000400C0060000040088323044201C850020820400101880",
INIT_05 => X"0200020040048A09202420000C00410402000025000800020804207000100800",
INIT_06 => X"10488704884D080202086A0A3429004012120004DC08125400A0008300821000",
INIT_07 => X"000800002C30204084381000128104000100002040003164040D800000400009",
INIT_08 => X"0440050003080202202400100080000000000C3E0408104C8000102300008810",
INIT_09 => X"4810240104111104200080120210A5104000A204615201500801010000AA10C0",
INIT_0A => X"81F525A82804010009029290200008B202238008080240000040100242048025",
INIT_0B => X"00A1141002C91844522A0004120488000800028000044000080020AF09240010",
INIT_0C => X"0408104081000810408100081040810008104040800408208040000008010121",
INIT_0D => X"4201E0B4000803200C150108008490809A002192462424202200440404204041",
INIT_0E => X"0804100160006000120002120499020A04A14650A32851962965190014200240",
INIT_0F => X"000000000080A200100021000000014020080021000000014020000014260082",
INIT_10 => X"0000000000000340080028000000014020080028000000014020008000008000",
INIT_11 => X"008000008000000000000081500010000100800000000000008C100080000012",
INIT_12 => X"05D0000880000006800058000020000000000005000000000000000048100100",
INIT_13 => X"0000D02E8040200000003401F80004000000000040026000274000900000001A",
INIT_14 => X"800023B8000030000000000042A00009AB00008800000000008012BA01001000",
INIT_15 => X"00A000106520350000040100000000000010C0200009BA000200000000000105",
INIT_16 => X"465196651B328CA8D26540544924272EB91004002022024048400000098030A0",
INIT_17 => X"6509425094250942509425094250942509425094250942509425094251946519",
INIT_18 => X"5094250942509425094250942519465194651946519465194651946519465194",
INIT_19 => X"2A05404808000000000000000014651946519465194651946519465094250942",
INIT_1A => X"69A69A69A68945B080201C92410480ABD102E689999E91BCD151200C30AE1C71",
INIT_1B => X"341A0D068341A0D068341A28A28A28A28A28A28A28A28A28A28A28A28A28A69A",
INIT_1C => X"FFC5B52068349A4D068341A0D269341A0D269341A0D068349A4D068349A4D068",
INIT_1D => X"0F7D17FFFFAAAE800000000000000000000000000000000000000000000003FF",
INIT_1E => X"EFAA843DE00F7803FEBAFFFFC2000557FEABEFA2D1400AA5D2AAAA00F7FFEAA1",
INIT_1F => X"4105555421EFF78028BEF5D003DFEFF7FFE8ABAF7802ABEFAAAE820000000021",
INIT_20 => X"AB45557BC0155007FFDEBAAA843DE00557BEAABAA2AEAABEFF78015555AA8017",
INIT_21 => X"154AAA2AA955FF00043DE005504175FF0851401455555555EFA2FBC01FFF7AAA",
INIT_22 => X"57DE105D2EBDF55557FFDE00552A974AAA2843DEAA5D2A820BA000428AAAAA84",
INIT_23 => X"517FFEFAAAEBDF45FFAEA8ABAF7D1400BAAAAE821EFF7D17DEAA5D2AAAAAA5D5",
INIT_24 => X"0000000000002ABFFA280154BAFF803DF45FFD17DFFFFFD56AA00557FC201000",
INIT_25 => X"4120ADA38E3F1EFA28F7DF7DFD7A2A4800000000000000000000000000000000",
INIT_26 => X"7A2A482038000A001C7A2803AE38FF843DEBAEBFFC20285D75EFBC7A2DB40082",
INIT_27 => X"C7EB8417555AA84104385D55421C7FF8028BEF41003FFD7F7F1EDA82F78E2DBD",
INIT_28 => X"5C7A2FBC51EFEBA0A8B6D5571C716D1475FFEAAA28E3FE385D71E8AAAAAA0A8B",
INIT_29 => X"50AA1C0428ABAB68E124BAA2AA955C708003FE285D00155FF0055451555D5F57",
INIT_2A => X"7FE825520ADA92495B7AE10412EBFF45497FFFE105D2E97482AA8038EAA412E8",
INIT_2B => X"F6DA284175C001000557FFEFB6A0BFF55F7AEAAA82FFDF40092B6A4871EFFFD5",
INIT_2C => X"0000000000000000000000000000028BEFA28E124AAF7843AF7DEBDB78FFFE3D",
INIT_2D => X"5517DF55A2FBC201008003DEAAA2D57FEAAF7FBFDF45AA800000000000000000",
INIT_2E => X"FFD57FE00FFAABFF45AA80020BA082E82155AA802AAAAFF803DEBAAAFBC20BA5",
INIT_2F => X"A5D5568ABAA2842AB55A28015545A284000BA5D5340145F78028BFF08003DF45",
INIT_30 => X"EF0855575455D7BD5555A2FBD75FFA2842ABFF5555575FF55557FEAAA2AABFEA",
INIT_31 => X"400A2802AABA002A954AA5D0028ABAF7AA820BAAAAE9754500043DEBA5D04175",
INIT_32 => X"2010FF80155EFF7D57DE005D003DE00007FEAA10002ABFF450079FFE005D2A97",
INIT_33 => X"2ABEFAAFFEABEFAAFFFDEAA00514200008517DFEFFF803FF45FFAAA8A00F7FBC",
INIT_34 => X"000000000000000000000000000000000000000000000028BFFA2AE820AAFF80",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000002000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033022000000180006",
INIT_01 => X"0000098218302849180060000C00424040000000080000080200090008510200",
INIT_02 => X"0801080200100000044008000080000041000000002002400800000009008010",
INIT_03 => X"0001000004000040000202000000000803006400088000003080040008C10000",
INIT_04 => X"0000100022008000000C08C00C00000400201830040000040000000400001820",
INIT_05 => X"0200000040000000248080210044000400000000000800000004000010000800",
INIT_06 => X"100007000049000202086A080000004010100000880800001000000030829000",
INIT_07 => X"000800002420000004201000128100000300002040003124040D802040400009",
INIT_08 => X"040005000108020220240020008000000000043E000000488000000100008811",
INIT_09 => X"0810040105111000202000024010A51040088080000000110000002000020084",
INIT_0A => X"040000000000010000040010200008B202230480080002000000100240008021",
INIT_0B => X"40003C020AC04400022808001000014000040088140000000000828000000820",
INIT_0C => X"0040004400044000040000400044000440000400002000221048840009012124",
INIT_0D => X"0002A00800000100440000000800800018002000008000800040022000000400",
INIT_0E => X"0804100100002000100002001001024800020001000080004000000800904000",
INIT_0F => X"000000000000A000102008000000014000082008000000014000000000240082",
INIT_10 => X"0000000000000240082001000000014000082001000000014000028000000000",
INIT_11 => X"028000000000000000000001400012000200000000000000000C100084000800",
INIT_12 => X"0000080000000004800000400020400000010000000000000000000048000000",
INIT_13 => X"0000900000010000000024080000000000000000000250002000200000000012",
INIT_14 => X"4000200000400000000000000290000100002000000000000000120000010000",
INIT_15 => X"0000001000000000010000000000000000104010000100000000000000000005",
INIT_16 => X"0000000001400080002100544924002A000004000020000080000000010032A0",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100400000000",
INIT_18 => X"0000000000000000000000000010040100401004010040100401004010040100",
INIT_19 => X"02A1410808000000000000000000000000000000000000000000000000000000",
INIT_1A => X"145145145146AB2A0CCC2A28A28A7AA0CDF0D1215281FC1A72E24C28E921AAA9",
INIT_1B => X"CA6532994CA6532994CA65145145145145145145145145145145145145145145",
INIT_1C => X"FFD9C63B95CA6532994CA6532B95CAE572994CA6532994CAE572B95CA6532994",
INIT_1D => X"FAAD1555FFF78400000000000000000000000000000000000000000000000200",
INIT_1E => X"AA5D2AAAA00F7FFEAA10F7D17FFFFAAAE801FF08557DF4555516AA00007BEABE",
INIT_1F => X"000557FC0010AAD57FF45A2D56AA0000043FFEFA2FFFDE1008556ABEFA2D1400",
INIT_20 => X"DEAA007FEAB45AAAE800AAF784020000000021EFAA843DE00F7803FEBAFFFFC2",
INIT_21 => X"421EFF78028BEF5D003DFEFF7FFE8ABAF7802ABEFAAAEA8BFF5D0415400F7FBF",
INIT_22 => X"015555AA80174105555401FF5D0415555557BFDFEF00517DE00A28028B450855",
INIT_23 => X"FFD7555AAD56AB45A2AE800AA5D7FFDEBAF7AEBDE00557BEAABAA2AEAABEFF78",
INIT_24 => X"000000000000155EFA2FBC01FFF7AAAAB45557BC0155007FFDEBAAA8417410AA",
INIT_25 => X"55556AA381C75EABEFBED1575C7E380000000000000000000000000000000000",
INIT_26 => X"81C516FBC7A2DB400824120ADA38E3F1EFA28F7DF7DFD7A2A4801EF085F7AF6D",
INIT_27 => X"38FF843DEBAEBFFC20285D75C0010AADF7AF6DB6D56FA3814003AFFFA2F1F8E3",
INIT_28 => X"BEF550412428F7F5FDE920875E8B45BEA0850BAE38002038000A001C7A2803AE",
INIT_29 => X"8E10AA802FB450851421C7FF8028BEF41003FFD7F7F1EDA82F78E2DBD7A2A4AD",
INIT_2A => X"E8AAAAAA0A8BC7EB8417555AA84104385D55401C75504125455575FAFD714557",
INIT_2B => X"5FFEAAA28E10438AAF5D2545BED56FB45BEA082082557BF8EBAF7AABFE385D71",
INIT_2C => X"00000000000000000000000000000175C7A2FBC51EFEBA0A8B6D5571C716D147",
INIT_2D => X"A80021FF007BE8BFF5D516AABA5D5568BEFF7D157555AA800000000000000000",
INIT_2E => X"5D002ABFFA2D16AAAA55517DF55A2FBC201008003DEAAA2D57FEAAF7FBFDF45A",
INIT_2F => X"A082E82155AA802AAAAFF803DEBAAAFBC20BA555140010AAFFE8BFFFFD17DEBA",
INIT_30 => X"00FFAABFF45AA803FFEF5500020BAFFD17DE10005568B55FF80154BAA280020B",
INIT_31 => X"1555D556AB555D5568A00AA843FF55085140145F78028BFF08003DF45FFD57FE",
INIT_32 => X"AAAAF7AABFEAA5D5568ABAA2842AB55A28015545A284000BA5D5342145550402",
INIT_33 => X"2ABFF5555575FF55557FEAAA2AA800AAAAD142155F7D57DF45FF8002010557FE",
INIT_34 => X"000000000000000000000000000000000000000000000015555A2FBD75FFA284",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000023FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B830084C1820E0000C36424840000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"000406A492E6E440842254D002108153422004800880000030C0315688C00006",
INIT_04 => X"00001201200090001205400000000094108C322644240C840008030440111800",
INIT_05 => X"222000444008010028404002A002009402400025080880000C04223000170900",
INIT_06 => X"12801628014B0B000A086CA6556800C012121004540816544522008200821100",
INIT_07 => X"1C08320054B624408428100094ADD080011721A04000316C140CA1A8A1F90019",
INIT_08 => X"00140500090B02C2E0EC04D1C08000000000647E858A104C920C81A5011088A6",
INIT_09 => X"40002481041F165820000101024061004004800567603592A801014C46426011",
INIT_0A => X"8404002020000101B0070310200008B60A23A51B28024CE24E40100260040004",
INIT_0B => X"2800340208811865D22BB384100E01090805A495100400050800E24D49A424C5",
INIT_0C => X"0C72A0872A0C72A0872A0C72A0C72A0872A0C595043950421400800009010104",
INIT_0D => X"4290A088812203360410110A400085539800210404C048CAC040464D28014405",
INIT_0E => X"0804101160006000101004A01811064B050204810240812241280D00200A0804",
INIT_0F => X"6D0141B0482A01AAEC3602330CD2A02952DC3502330CB4A0318B414000240082",
INIT_10 => X"5B4551630144C0155C3502330CD2A02952DC3602330CB4A0318B5600C587149B",
INIT_11 => X"FE04E587083B6A51005956308D1E8202C436375908AA840AD4513437640F1524",
INIT_12 => X"E020C67062F47B2872400044959BC42B1060F0D036B80B548523136C158878D8",
INIT_13 => X"8F0B27010A2699AAA3794392000D81852B0A050C224180062085134CD1719564",
INIT_14 => X"0AD57400C50500D94C8121713C02B555101C90705D71009604140C0418CE0C37",
INIT_15 => X"DC06A27C828E024D8C50965A40821568A06113801505010334AA73AA0666DAC2",
INIT_16 => X"04812048123408C0822040004C248604B2100400100084008001D0113920060C",
INIT_17 => X"4812048120481204812048120481204812048120481204812048120481204812",
INIT_18 => X"8020080200802008020080200812048120481204812048120481204812048120",
INIT_19 => X"00A0014200000000000000000020080200802008020080200802008020080200",
INIT_1A => X"4104104104140D220A4A380000002A80E900C4C1100830181621409C80210821",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000410",
INIT_1C => X"FFC1F83800000000000008040000000000000000000201000000000000000000",
INIT_1D => X"0F7842AA00002A80000000000000000000000000000000000000000000000200",
INIT_1E => X"4555516AA00007BEABEFAAD1555FFF784020AAF7D542155F7D1400AAF7FFFDE0",
INIT_1F => X"FFFAAAEA8ABAFFD17FEBAFFAA800AA007FFDFFFA28428A000000001FF08557DF",
INIT_20 => X"00AAF78028AAAFF84020AAFFFBEABEFA2D1400AA5D2AAAA00F7FFEAA10F7D17F",
INIT_21 => X"40010AAD57FF45A2D56AA0000043FFEFA2FFFDE1008556AB45555568A10A2FFC",
INIT_22 => X"03FEBAFFFFC2000557FC0155FFD1555FF0804000AA000428A10AAAA801EFFFD1",
INIT_23 => X"8428A10087FD7400552EBDFEFA2FBFFF550000020000000021EFAA843DE00F78",
INIT_24 => X"00000000000028BFF5D0415400F7FBFDEAA007FEAB45AAAE800AAF78428B45A2",
INIT_25 => X"E3DF450AAF7F1FDE38FF8A2DA101C2A800000000000000000000000000000000",
INIT_26 => X"01C0E001EF085F7AF6D55556AA381C75EABEFBED1575C7E380000BAF7DB4016D",
INIT_27 => X"38E3F1EFA28F7DF7DFD7A2A4AFABAFFDF7AE82F7AA870AA0071F8FFFBE842DA1",
INIT_28 => X"B455D5B68A28A2FFC20AAEB842DAAAE38A02082E3FBEFBC7A2DB400824120ADA",
INIT_29 => X"8A28AAA4801FFE3DF40010AADF7AF6DB6D56FA3814003AFFFA2F1F8E381C516D",
INIT_2A => X"001C7A2803AE38FF843DEBAEBFFC20285D75C2145F7DF525EF140A050AA1C002",
INIT_2B => X"0850BAE3802DB6DAA8A28A00007FD74284120BFFFFBEF1F8F7D080A02038000A",
INIT_2C => X"000000000000000000000000000002DBEF550412428F7F5FDE920875E8B45BEA",
INIT_2D => X"A80020BAFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE10552E8000000000000000",
INIT_2E => X"085568BEFF7803FE10552E821FF007BE8BFF5D516AABA5D5568BEFF7D157555A",
INIT_2F => X"5A2FBC201008003DEAAA2D57FEAAF7FBFDF45AA803FEBAFFFBEAA00F7AE974BA",
INIT_30 => X"FFA2D16AAAA55517DF55557FEAAAAA2FFC00AAAA803FEAAA2AA82000A2FFFDF5",
INIT_31 => X"1EF552E974BA550028ABAA280001FFAAFFC0010AAFFE8BFFFFD17DEBA5D002AB",
INIT_32 => X"ABFF082E820BA082E82155AA802AAAAFF803DEBAAAFBC20BA555142155F7FFC0",
INIT_33 => X"7DE10005568B55FF80154BAA2803FFFFA2AAAAA00007FD74BA08003DFFFFFD16",
INIT_34 => X"00000000000000000000000000000000000000000000003FFEF5500020BAFFD1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000002000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C048000C048400380000007026040000000080000088200002802153231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"210D050012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"0080100022408000060DE0000066630C70241827041000040800820480001AA4",
INIT_05 => X"0240000C400000003C808003E0C8001401000000040900020904004000070800",
INIT_06 => X"1800068000491300CF0969A421C0004018184000100804005784000130821200",
INIT_07 => X"7E8C53200CA4850224301807D1CB45900147E03040083124FC0CD0C8A1FF0019",
INIT_08 => X"0046050013081206A4A503A9E8C0812000001C7E11A24058B84D40E33992D98F",
INIT_09 => X"010004810491175C20000080000821004010C01086003C13E000004EDF020400",
INIT_0A => X"000000000000010000180018200408B27E234913E9000CFA09A8180248001000",
INIT_0B => X"ACA0141000800021826933E03662802B3001E09F000000023000000000000867",
INIT_0C => X"0832F0C32F0832F0832F0C32F0832F0832F0C197861978400000000208010100",
INIT_0D => X"05FA0201E7F3F01F40401C17E800C7F3380020000000006AE01180493C5BC1AF",
INIT_0E => X"000200F500002200004005002001408400000000000000000000053A4096F807",
INIT_0F => X"246FC1B17B2C53F2FC16691DB587201EDDF4162B1DB527201EDDC46070241001",
INIT_10 => X"2A67DF2A01D5CC9794162B1DB587201EDDF416691DB527201EDDD884272592D6",
INIT_11 => X"288007258E995D5A825DBA569F9FF02547068618CD3CC45B7863AE7EC00D4B12",
INIT_12 => X"F6208C6CCA5C33717461C045B5B182019473D19D7CCD856106F31A683621BDFC",
INIT_13 => X"866E2FB10A652CC8E3538BBA01624E51AA6C0469AC5493F5688532966471A9C5",
INIT_14 => X"4F9B740041E1F5759001B4AA1853E6D5144AA9C914C8608D2724A4C4118D992B",
INIT_15 => X"DE07EAD9825682D4A36C0B0B4B85112B2C4A05D3E6D5051893335EB0072AA85A",
INIT_16 => X"00000000008000000821000048260020000004001DC0800000010E7F70171401",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0100401004010040100401004000000000000000000000000000000000000000",
INIT_19 => X"2A21010808000000000000000000401004010040100401004010040100401004",
INIT_1A => X"4924924924890380800016A28A28802B10B83728C1111026C152A23010848658",
INIT_1B => X"6432190C86432190C86432082082082082082082082082082082082082082492",
INIT_1C => X"FFDE003AC964B2592C964B2592C964B2592C964B2592C964B2592C964B2592C9",
INIT_1D => X"5FFAA80155F78400000000000000000000000000000000000000000000000200",
INIT_1E => X"55F7D1400AAF7FFFDE00F7842AA00002AAAA10FF8002155F7FFC200008041755",
INIT_1F => X"5FFF7842AB55080000145557FE8AAA080000155F7FFFDEAA0000020AAF7D5421",
INIT_20 => X"2000FF80020AAA2AAAABFF002E801FF08557DF4555516AA00007BEABEFAAD155",
INIT_21 => X"A8ABAFFD17FEBAFFAA800AA007FFDFFFA28428A00000028B4555043DFFFFFAE8",
INIT_22 => X"FEAA10F7D17FFFFAAAE80000A284174AAFF8428AAAFF8415545AAFBD7545F7AA",
INIT_23 => X"00000105D55400AA082A82155F7FFFDEAA08556ABEFA2D1400AA5D2AAAA00F7F",
INIT_24 => X"0000000000002AB45555568A10A2FFC00AAF78028AAAFF84020AAFFFBC215508",
INIT_25 => X"E3F5C000014041256DEBA487145F784000000000000000000000000000000000",
INIT_26 => X"2080E000BAF7DB4016DE3DF450AAF7F1FDE38FF8A2DA101C2AAFA00EB8E0516D",
INIT_27 => X"381C75EABEFBED1575C7E3802FB551C0E0516D417FEDA921C000017DEBF5FDE9",
INIT_28 => X"B55410A3FFC7F7A087000FF80070BAAAAAADBD70820801EF085F7AF6D55556AA",
INIT_29 => X"556DA2FBD7545F7AAAFABAFFDF7AE82F7AA870AA0071F8FFFBE842DA101C0E2D",
INIT_2A => X"400824120ADA38E3F1EFA28F7DF7DFD7A2A480000BE8A17482F78A28A92E3841",
INIT_2B => X"A02082E3FBC217D1C0E0500041554508208208017DF7F5FDE9208556FBC7A2DB",
INIT_2C => X"000000000000000000000000000002DB455D5B68A28A2FFC20AAEB842DAAAE38",
INIT_2D => X"52EBDE00AAAE975FFAAD1420005504001FFAA8015545F7800000000000000000",
INIT_2E => X"5504001FFAAD17DE00082E820BAFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE105",
INIT_2F => X"F007BE8BFF5D516AABA5D5568BEFF7D157555AA803DF45552E975EF007FFFE00",
INIT_30 => X"EFF7803FE10552EBDF45002EBFF55FF8017410FF84154BAAAAABFF450000021F",
INIT_31 => X"400F7AEA8A10A284175FFAAFBD5555F7AEBFEBAFFFBEAA00F7AE974BA085568B",
INIT_32 => X"DE1008517DF55A2FBC201008003DEAAA2D57FEAAF7FBFDF45AA8002000FFAE95",
INIT_33 => X"C00AAAA803FEAAA2AA82000A2FFC21EF552A954100851554000004021FFFFD17",
INIT_34 => X"00000000000000000000000000000000000000000000003DF55557FEAAAAA2FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00010100926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"0004122122029100100C00001200009C40A83A2044360C84190BAC04E0101820",
INIT_05 => X"027000004009050064C8C00104C10184034010250089C00EB004327064B60900",
INIT_06 => X"1B9416B94149000402086D42142800C012125804440812541027008230821380",
INIT_07 => X"0008320014B02848A4A8100015C55500057801A04000712C040CB1F880600009",
INIT_08 => X"005005000908020220E40170008042000000557E048A144C800590010000882D",
INIT_09 => X"0100250104B5310020000100020821004016CC1C616401910801010100CA2040",
INIT_0A => X"800000000000010192072310200028B6022346080802C0074AC0100259001004",
INIT_0B => X"A8201410008088C5D2288004120E802908800488000500050800404D49A42EB0",
INIT_0C => X"0400000000040000000000000040000000000000020000000000000008010102",
INIT_0D => X"4A02008000000360401021280800E400B800610C844848200028448400000000",
INIT_0E => X"000000086000600040D045E4195104D5854284A14250A12A512A880828984008",
INIT_0F => X"85D480949E07A80948354B6E68982167061037496E6838216706206810240000",
INIT_10 => X"652138E510B456587037496E689821670610354B6E6838216706220431961CA9",
INIT_11 => X"C2043196186A91674011CE61403562274AA49CD594CF00039C7C414B6509DA22",
INIT_12 => X"8A2E6A983014780CC8604040424A5323845932E620295879818170304B2F5002",
INIT_13 => X"8F019451654B9104A328665603148895D44E0251142B42A3D8B2A5C882519432",
INIT_14 => X"0AC5DC06A6C6A465AA0091482382B17614F2202858EE300991415B45CD530602",
INIT_15 => X"4000052E08DC8047F17D1C7C3C02128E587D6A02B17605A130A4E8BF00225885",
INIT_16 => X"84A1284A123508508220808048240604B2100C00022084809000D000393722A1",
INIT_17 => X"4A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A12",
INIT_18 => X"A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A128",
INIT_19 => X"F1228154000000000000000000284A1284A1284A1284A1284A1284A1284A1284",
INIT_1A => X"75D75D75D75FFAFEFEFEEEAAAAAAFBF3FC1FF77DDFE7EFBEFFE7CFC0044FBEFB",
INIT_1B => X"FAFD7EBF5FAFD7EBF5FAFD75D75D75D75D75D75D75D75D75D75D75D75D75D75D",
INIT_1C => X"FFC0003BF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5",
INIT_1D => X"F007FE8A00AAFBC0000000000000000000000000000000000000000000000200",
INIT_1E => X"55F7FFC2000080417555FFAA80155F7842AB55552E821FFFFD5555EF552ABDFE",
INIT_1F => X"A00002A821EF5D7BC21FFFFFBD55EFAAD1554BA00556AA00AAD16AA10FF80021",
INIT_20 => X"FF45A2AABFEBA082A975555D55420AAF7D542155F7D1400AAF7FFFDE00F7842A",
INIT_21 => X"EAB55080000145557FE8AAA080000155F7FFFDEAA00002AB45082A821EF5D557",
INIT_22 => X"BEABEFAAD1555FFF7842AABAA2FFE8BEF5D517FF455D554214500043DEBAAAFF",
INIT_23 => X"AABDF555D2E955EFA28428A10552EBFEAAAAD1401FF08557DF4555516AA00007",
INIT_24 => X"00000000000028B4555043DFFFFFAE82000FF80020AAA2AAAABFF002E80000AA",
INIT_25 => X"EBD5525C74124B8FC71C71EFA28AAF5C00000000000000000000000000000000",
INIT_26 => X"8AAD16FA00EB8E0516DE3F5C000014041256DEBA487145F78428B6D4120851FF",
INIT_27 => X"AAF7F1FDE38FF8A2DA101C2A871C74975C01FFEBF5D25EFA2D555482085F6FA2",
INIT_28 => X"B7D1C24851FF495F7FF55A2A0BFE921C2E9557D415B400BAF7DB4016DE3DF450",
INIT_29 => X"214508003FEAABEFFEFB551C0E0516D417FEDA921C000017DEBF5FDE92080E2A",
INIT_2A => X"7AF6D55556AA381C75EABEFBED1575C7E38028A82B6F1E8BFF495F78F7D49554",
INIT_2B => X"AADBD7082087000AAA4BFF7D5D20905C7AA842DA00492EBFEAABED1401EF085F",
INIT_2C => X"000000000000000000000000000002DB55410A3FFC7F7A087000FF80070BAAAA",
INIT_2D => X"78028BFF0004175EFA2D54214508042AB455D517DEBAA2D54000000000000000",
INIT_2E => X"AAD557410007BFDEAAA2D57DE00AAAE975FFAAD1420005504001FFAA8015545F",
INIT_2F => X"AFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE10552E975450051401EFA2D5421EF",
INIT_30 => X"FFAAD17DE00082EA8BFF5504175FF087BFFF45AA843FE005D2A955FF087BC20B",
INIT_31 => X"BFF087BEABEF00554215500003FEBAFFFBFDF45552E975EF007FFFE005504001",
INIT_32 => X"FEAAFFD5421FF007BE8BFF5D516AABA5D5568BEFF7D157555AA8028A00FFD16A",
INIT_33 => X"17410FF84154BAAAAABFF45000017410AA803DFEF550402155A2843FE00082AB",
INIT_34 => X"00000000000000000000000000000000000000000000003DF45002EBFF55FF80",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000033FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"000103A7A00904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000120122009000100C00000000000400A83A2044200C840000800400101820",
INIT_05 => X"020000004008010024C0C0010040000402000025000800020004207000100800",
INIT_06 => X"108016080149080002086807542800C012120004440812541020008230821000",
INIT_07 => X"4008120054B42850B42A100010ED1500010001A040003164040CF5E201400009",
INIT_08 => X"00400500090A020220A40A7000800000000014FE8508144C924080C100008801",
INIT_09 => X"0000040104111100200001000200210040008004616001910801010000422000",
INIT_0A => X"800000000000010190070310200008B202236D080802400002C0100240000000",
INIT_0B => X"0000141000800844522800041204000008000488000400000800004D49240820",
INIT_0C => X"0400004000000000000004000000000000004000000000000000000008010100",
INIT_0D => X"42020080000002204010010808008000B8002104044048200000440400000000",
INIT_0E => X"0000000000006000000000201811004005020481024081224128080820984000",
INIT_0F => X"CBA340480040A100A42008000161C140000420080001C1C14000032010240000",
INIT_10 => X"1A8A039600022260042001000161C140000420010001C1C140001604E8084341",
INIT_11 => X"1E04E8082580E2B8802201014800C220A21829A302F1C024010C001124020C8C",
INIT_12 => X"0024ACA60CA000048228404401004418012787124648157780120B8678C00080",
INIT_13 => X"00009001072D04730000241000CB1325E78E0186030240000083B60239800012",
INIT_14 => X"00001001EF6F4163C480481506800004000CFD55196CB012481812049495C194",
INIT_15 => X"40068248800108B8FB61A0401200845594965000000400568D0CFB7800550605",
INIT_16 => X"04812048123408408220000048240604B210040000008400800B0000090022A1",
INIT_17 => X"4812048120481204812048120481204812048120481204812048120481204812",
INIT_18 => X"8120481204812048120481204812048120481204812048120481204812048120",
INIT_19 => X"2820014000000000000000000020481204812048120481204812048120481204",
INIT_1A => X"3CF3CF3CF3CFFBBEEEEEFE79E79EFAABDDFAF369CB91FE1EF7D3AEBBDBAFBEFB",
INIT_1B => X"FE7F3F9FCFE7F3F9FCFE7F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"FFDFFFC1FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"AAAAEAAB45082E80000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFD5555EF552ABDFEF007FE8A00AAFBE8BEFA2D568ABA00003DF555555574A",
INIT_1F => X"155F78428AAA007FE8A1008002AABA555155400557BC2010557BEAB55552E821",
INIT_20 => X"FFFF082EBDEBAA2D1420105D002AA10FF8002155F7FFC2000080417555FFAA80",
INIT_21 => X"C21EF5D7BC21FFFFFBD55EFAAD1554BA00556AA00AAD140145AA8028ABA002EB",
INIT_22 => X"FFDE00F7842AA00002A80155A2AEA8A10080428A10FFAEBFFEF5D0428B45A2FF",
INIT_23 => X"5568A000000175FFF7D155545F7FBC0010FFAA820AAF7D542155F7D1400AAF7F",
INIT_24 => X"0000000000002AB45082A821EF5D557FF45A2AABFEBA082A975555D55400BA00",
INIT_25 => X"000E38F6D4155504AAA2AEAAB6D0024800000000000000000000000000000000",
INIT_26 => X"05D75E8B6D4120851FFEBD5525C74124B8FC71C71EFA28AAF5E8BFFB6D56DA82",
INIT_27 => X"0014041256DEBA487145F78428ABA147FEDA10080E2AAAA555552400417FC200",
INIT_28 => X"155BE8028A82002EB8FC70024BAEAAB6DB4202849042FA00EB8E0516DE3F5C00",
INIT_29 => X"DFD7550428B55A2F1C71C74975C01FFEBF5D25EFA2D555482085F6FA28AAD147",
INIT_2A => X"4016DE3DF450AAF7F1FDE38FF8A2DA101C2A80145B6AEA8A10080E2DA00F7A0B",
INIT_2B => X"E9557D415B400AA00556DA000004175FFE3D15757DE3F5C0038FFAA800BAF7DB",
INIT_2C => X"000000000000000000000000000002AB7D1C24851FF495F7FF55A2A0BFE921C2",
INIT_2D => X"2D568BEFFFD57FE10002AAABEF0051400AAA2AAAABFF08000000000000000000",
INIT_2E => X"5D5142000007BC20105D5568BFF0004175EFA2D54214508042AB455D517DEBAA",
INIT_2F => X"0AAAE975FFAAD1420005504001FFAA8015545F78028AAA557FFFE00082EAAAAA",
INIT_30 => X"10007BFDEAAA2D557555FF8028A00082EAAB45000028ABAFFFBC20AA08043DE0",
INIT_31 => X"A10002ABFE00F7803FF555D002AB55AAD1575450051401EFA2D5421EFAAD5574",
INIT_32 => X"20BAFFAE820BAFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE10552E82155FFAAA8",
INIT_33 => X"FFF45AA843FE005D2A955FF087BC20AA00517DE000804175EFAAD1555EFA2D14",
INIT_34 => X"000000000000000000000000000000000000000000000028BFF5504175FF087B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000080000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"0001100024A0800000440000000000040088322044200C840000011400151800",
INIT_05 => X"A200014C4000000020000000000B8094020000254C8800000514203000108800",
INIT_06 => X"10000600004B0044020868021428004012120005540812540020008600831000",
INIT_07 => X"00086100043224489428100010811100010001A040003124040CAC6000400009",
INIT_08 => X"00160500090A0282A06400100080C300000005BE0488104C8000000100008800",
INIT_09 => X"00000581041110022000000002002100400080046140011008010100008A0400",
INIT_0A => X"800000000000010180060210200008B2022304080800400007C0100240000000",
INIT_0B => X"0004140000800844522800041004000008000080000400000800000D09240000",
INIT_0C => X"0400004000040000400000000000000000004000020000200000000008010100",
INIT_0D => X"4A00008000000260001001280000C400B0002000000000000000440400000000",
INIT_0E => X"0000000840006000000000001001004004000000000000020100000000000000",
INIT_0F => X"0000000000000000002021000000000000002021000000000000046000240000",
INIT_10 => X"0000000000000000002028000000000000002028000000000000020000008000",
INIT_11 => X"0200000080000000000000000000020001008000000000000000000004000012",
INIT_12 => X"0020000880000000006000400080C0000000000D081202800000000000000000",
INIT_13 => X"0000000100402000000000100000040200100000000000000080009000000000",
INIT_14 => X"0000100000003088014000000000000400000088221100000000000401001000",
INIT_15 => X"4000000800000000048407170500000000000000000400000200000000000000",
INIT_16 => X"00000000023000000220000048240404A010040000008000000000000000020C",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0020014000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000020000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFC0000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"555003DE10A2FBC0000000000000000000000000000000000000000000000200",
INIT_1E => X"BA00003DF555555574AAAAAEAAB45082EBFE000004020AA552E80000F7FBC214",
INIT_1F => X"A00AAFBFDEBA555568BEFA2FBE8A10F7802AA0055003FE10007BE8BEFA2D568A",
INIT_20 => X"55EFF78428BEFAAD17DF55AAAEAAB55552E821FFFFD5555EF552ABDFEF007FE8",
INIT_21 => X"28AAA007FE8A1008002AABA555155400557BC2010557BFFFEFA2FFC20005D2A9",
INIT_22 => X"417555FFAA80155F7843DF455D2AA8B45AAD57FF55A2FBC21FFA28415400FF80",
INIT_23 => X"514200055002AA00AA802AABA002E9740055516AA10FF8002155F7FFC2000080",
INIT_24 => X"00000000000000145AA8028ABA002EBFFFF082EBDEBAA2D1420105D003FFFF08",
INIT_25 => X"412A87010E3F5C0145410E3DE28B6FFC00000000000000000000000000000000",
INIT_26 => X"8147FE8BFFB6D56DA82000E38F6D4155504AAA2AEAAB6D0024B8E381C0A00092",
INIT_27 => X"C74124B8FC71C71EFA28AAF5F8EAA495F68BFFA2F1EFA38E38428A005D0038E2",
INIT_28 => X"FFFBEF5C0000492A955FFF78428BEFB6DB7DF45AAAEA8B6D4120851FFEBD5525",
INIT_29 => X"21EFAA8E10400E38E28ABA147FEDA10080E2AAAA555552400417FC20005D75F8",
INIT_2A => X"0516DE3F5C000014041256DEBA487145F7843FF7D4120A8B6DAAD17FF55B6F5C",
INIT_2B => X"B4202849043FFC7005F4501041002FA38A2842AA82142095428415F6FA00EB8E",
INIT_2C => X"0000000000000000000000000000007155BE8028A82002EB8FC70024BAEAAB6D",
INIT_2D => X"8002AAAA5D2A82000082E95400A2D542155002ABDEBAF7FBC000000000000000",
INIT_2E => X"A2802AA105D002AABA5D7BE8BEFFFD57FE10002AAABEF0051400AAA2AAAABFF0",
INIT_2F => X"F0004175EFA2D54214508042AB455D517DEBAA2D56AABA087BEABEFAAD57DEAA",
INIT_30 => X"00007BC20105D556ABFFF7D142010082A955EFFF8428BFFFFFBFDF55A2AEA8BF",
INIT_31 => X"BEFA2D57DF45F7D1401FFA2AA82000AAAAA8AAA557FFFE00082EAAAAA5D51420",
INIT_32 => X"54AA007BFDE00AAAE975FFAAD1420005504001FFAA8015545F7803FFEF08002A",
INIT_33 => X"AAB45000028ABAFFFBC20AA08043FF55087BD740000043DEAAA2842AA005D001",
INIT_34 => X"000000000000000000000000000000000000000000000017555FF8028A00082E",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000003000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"010108A802BB00080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"8BFA58800005C40A46240252145148B38248030356415A4E62B6FC660F287240",
INIT_05 => X"0F05EA11E570000D610000000710296E542B6E3A825C15FB30A643695BFC2D56",
INIT_06 => X"00000200021100C87570B08224C8AB52C0A8030140BCC0460050690A95C8383D",
INIT_07 => X"76F500240510A00205F0A407D0021A155378900002A002433A0AA00EE6E79564",
INIT_08 => X"00015995440C8327241440096A2800002828123D542910380004E03103624040",
INIT_09 => X"0010222D90409A05B2CB2CA400200209E5601044A24000000462A60018880100",
INIT_0A => X"300000000000259200140001A15000017F0051D0F837248C005514AC40C08205",
INIT_0B => X"395012004240014891801000495D40192D100000000005452D54000C09070003",
INIT_0C => X"6110001100011000110001100011000110001080008800080005202280801080",
INIT_0D => X"BB4000140A80A5C8000102ED0044008004AD324000000008003561180063DB4F",
INIT_0E => X"1400404912AA28AA890BA00000024800480000000000000200802151025062C0",
INIT_0F => X"6D0031F554E11C596A64003195933741477264003195555B418687E358360208",
INIT_10 => X"41CD50A499CF47DCB264003195933741597264003195555B4198843940076D29",
INIT_11 => X"043D400758486A556489347FE5F409CBC1362510695B6288743123C952518520",
INIT_12 => X"B1C74424EAE2992046EB70026486035600CEC45CBCA809654B48163CCC895E1E",
INIT_13 => X"C383298E3A242DEA151848302BFD6D522B10C7EC71F6C1DB071D1216E078C4C1",
INIT_14 => X"8B93D037DAAABC982BE22267A2E2E4F44AA1DC5E37400C9EE1B7B638E8849D23",
INIT_15 => X"86E6A2EE015998B28654565A003F0068E35352C1CAE48BFBF3A6C9B7B286B4DA",
INIT_16 => X"00000000009000040A8000452110A8442040D655602A102A0027E2C423202840",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"B020000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"28A28A28A28F4EF2FC3C34F3CF3C2AC31DF7A22A898D21B4C9838D30B6A7B451",
INIT_1B => X"F4FA3D3E8F4FA3D3E8F4FA68A68A68A68A68A68A68A68A68A68A68A68A68A28A",
INIT_1C => X"FFC00003E9F4FA7D3E9F47A3D1E8F47A3D1E8F47A3D3E9F4FA7D3E9F4FA7D3E9",
INIT_1D => X"AFF80001FF002A80000000000000000000000000000000000000000000000200",
INIT_1E => X"AA552E80000F7FBC214555003DE10A2FBC21FFFFFBFDF45A2D56AB45FFFFD54B",
INIT_1F => X"B45082E974BA5D7BFDF55A2FFFFE005D7BC0010002E954AA087FFFE000004020",
INIT_20 => X"7410FFD1555550000020BAAAFFE8BEFA2D568ABA00003DF555555574AAAAAEAA",
INIT_21 => X"BDEBA555568BEFA2FBE8A10F7802AA0055003FE10007BC0000082A9740055001",
INIT_22 => X"ABDFEF007FE8A00AAFBD55EFAAFBD74105504021FF5D2EAAABAFFFBD55FF002A",
INIT_23 => X"517DF45AAFFFFEAAFFAABFE10007FC00AA087FEAB55552E821FFFFD5555EF552",
INIT_24 => X"0000000000003FFEFA2FFC20005D2A955EFF78428BEFAAD17DF55AAAE820AA5D",
INIT_25 => X"AADB6FB6DFFFBD54AAE38E021FF0824800000000000000000000000000000000",
INIT_26 => X"A1C7FF8E381C0A00092412A87010E3F5C0145410E3DE28B6FFC21C7E3F1F8F55",
INIT_27 => X"6D4155504AAA2AEAAB6D002492482497BFDF45AAFFF8E385D7BC5000002E904B",
INIT_28 => X"010142E90428490015400FFDB555450804070BABEF5E8BFFB6D56DA82000E38F",
INIT_29 => X"DAAAFFF1D55FF002EB8EAA495F68BFFA2F1EFA38E38428A005D0038E28147FC2",
INIT_2A => X"851FFEBD5525C74124B8FC71C71EFA28AAF5D25D7B6F1D54384904021FF5D2AA",
INIT_2B => X"B7DF45AAAE820925D5B7DF45A2F1FDEAAEBAABDE001471C20921475E8B6D4120",
INIT_2C => X"0000000000000000000000000000038FFFBEF5C0000492A955FFF78428BEFB6D",
INIT_2D => X"7FBC2145AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF00000000000000000000",
INIT_2E => X"557FD7410082A800AA557BEAAAA5D2A82000082E95400A2D542155002ABDEBAF",
INIT_2F => X"FFFD57FE10002AAABEF0051400AAA2AAAABFF080000000087BFDF55A2FFE8AAA",
INIT_30 => X"105D002AABA5D7BC20005D2E800BA080417400F7FBD75450800174AAFFD168BE",
INIT_31 => X"4AA0800001EF5D2ABDEBAF7D1575EF082EAAABA087BEABEFAAD57DEAAA2802AA",
INIT_32 => X"0000555568BFF0004175EFA2D54214508042AB455D517DEBAA2D540155F7D155",
INIT_33 => X"955EFFF8428BFFFFFBFDF55A2AE82010557FFDF55A2D57FEAAAAAEBFE1055514",
INIT_34 => X"00000000000000000000000000000000000000000000002ABFFF7D142010082A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000001000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"294ADB4AFFCBF0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"DB7A40806FE4040840EBC563A0150A0926146FECB04196482236FC2005282AE1",
INIT_05 => X"0403DA0383200831C68206D7E6D0250834336D1E81500FDB306045255BFC2076",
INIT_06 => X"D0002200022D1C59E53558D3EBFC6701CBC303163670497AFF00291B3C0E2015",
INIT_07 => X"F81684248A38B022475DCA9BD00116E33CC3821774BB55F53BB42329AA3C0CEA",
INIT_08 => X"1660700CE0641527241060AD844E1C0088001223022D189A2800542219204903",
INIT_09 => X"B6D94C1C1C51DFF881861CBE0305A12A0321810217C01D34EDC98FFA1C8E0000",
INIT_0A => X"F1F1FD8F8FBDE40E001E000B3A5DAADAFDDA5DA79350DF70027CE86F047BEF19",
INIT_0B => X"2DD8141817C00319F8E853E64D73A08BFF00E9A7415606747E6610052CDEE97F",
INIT_0C => X"4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A7800617112E46F05D0",
INIT_0D => X"BFF252D4CFEB69FF7A5F5AFFCCA787F7FE67C2180000006CE8A3F06ABD73DBCF",
INIT_0E => X"94BB02C9F99FD0678B87A0003000D8D02E00000000000000040025D3C21463D6",
INIT_0F => X"6D2BF232221ABD9CA854DFDD64A67D42C0F054DFDD64667D42C063E57A8F7B45",
INIT_10 => X"EFBB5AEDAA504801F054DFDD64A67D42C0F054DFDD64667D42C07237DFE5865F",
INIT_11 => X"3A33DFE58EAE7F5AB50D0806A9A2E0DFFF47DEDC496DA3181A0CC71440F9FBC3",
INIT_12 => X"7056E9C9C3FC95949AEFF556EF9C75E7DCF1EB1B6E6FCDC87CB35FC94B36AECF",
INIT_13 => X"92B29382AF5B6AAAE594A4C0DBFDAD94AA669809809FEFAF4157ADB55572CA52",
INIT_14 => X"BEBF41AE33F32ADD543430808BABAF50E1A5EB4BAEA45A250202FE0ADD39387F",
INIT_15 => X"E83FB669523E865D4B1293AB6B90BF2F0E30EDEFAFD0B3FBD72E9E90D20A003F",
INIT_16 => X"0000000002F840000BCE0B6F67B3F845E017C833F6AAC02B002A2EFF22D4073D",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"CC0C006000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"34D34D34D352324C3434C0EBAEBA21BBE5F04006013DB9880A5D25C3230B88A7",
INIT_1B => X"1A0D06A351A0D06A351A0D34D75D34D34D75D34D75D34D34D75D34D75D34D34D",
INIT_1C => X"FFC00002351A8D46A351A8D46A351A8D46A351A8D468341A0D068341A0D06834",
INIT_1D => X"0007BEAB55FFAA800000000000000000000000000000000000000000000003FF",
INIT_1E => X"45A2D56AB45FFFFD54BAFF80001FF002A821FFFFFFFFFFFFFFBFDFEFAAD14201",
INIT_1F => X"E10A2FBEAB45A28000010082A975EFA2D140145007BC21FF5D2A821FFFFFBFDF",
INIT_20 => X"54AA0855575FFAAD57FE005D7BFFE000004020AA552E80000F7FBC214555003D",
INIT_21 => X"974BA5D7BFDF55A2FFFFE005D7BC0010002E954AA087FD7400082E954AA08001",
INIT_22 => X"5574AAAAAEAAB45082EBFFFFF7D16AB45FFFFEABEF007BD74005555555EFF7AE",
INIT_23 => X"84154BA082E801FFAAFBC0155555568B45552EA8BEFA2D568ABA00003DF55555",
INIT_24 => X"00000000000000000082A97400550017410FFD1555550000020BAAAFFC0145AA",
INIT_25 => X"F7F1FAFD7A2D5400001C7BEDB7DEBA4800000000000000000000000000000000",
INIT_26 => X"F4124821C7E3F1F8F55AADB6FB6DFFFBD54AAE38E021FF0824851FFFFFFFFFEF",
INIT_27 => X"10E3F5C0145410E3DE28B6FFEFB45AA8E070281C20925FFBEDB451451C7BC01E",
INIT_28 => X"4280024924AA1404174AA0055505EFBEDB7AE385D7FF8E381C0A00092412A870",
INIT_29 => X"54005D5B575EFEBAE92482497BFDF45AAFFF8E385D7BC5000002E904BA1C7FD5",
INIT_2A => X"6DA82000E38F6D4155504AAA2AEAAB6D0024BFFD7FFDB6AB7DFFF5EDBC71C7BD",
INIT_2B => X"4070BABEF5C516DAA8A124921C20801FFB6F5C0145555B68B7D4124A8BFFB6D5",
INIT_2C => X"0000000000000000000000000000002010142E90428490015400FFDB55545080",
INIT_2D => X"000155FFF7FBFDFEFFFD568B45AAD5400005D7BFFFEFAA800000000000000000",
INIT_2E => X"FFFFD5545557BC21FF080002145AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF0",
INIT_2F => X"A5D2A82000082E95400A2D542155002ABDEBAF7FBFDF55A2AA974AA5D04001EF",
INIT_30 => X"10082A800AA557BD74BA0004000AA5500174AA0855421FFFFFBEAAAA5D7BEAAA",
INIT_31 => X"BFFF7D57FF455D7FD54105D7BD75FFAAAA80000087BFDF55A2FFE8AAA557FD74",
INIT_32 => X"8BEF000028BEFFFD57FE10002AAABEF0051400AAA2AAAABFF08003FF55F7FFEA",
INIT_33 => X"17400F7FBD75450800174AAFFD1555FFA2AA800105504001EFFFD140145557BE",
INIT_34 => X"0000000000000000000000000000000000000000000000020005D2E800BA0804",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000033FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"0405D434003F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"50805AC31007D6125724029216554A9847669903D640EC8E2001002604503004",
INIT_05 => X"07008000E0EA11803850C800010022660C1C0065003C0404002646DC20A02D40",
INIT_06 => X"30A03A0A138900001127A09234C81FF040000000002C44D620F0228454C83810",
INIT_07 => X"405584280B10014003A8067400920810FF3C72024300A0030048221ACEE383E4",
INIT_08 => X"1000C983E6041505253500F66E620428000B1804000152E52801A20200840900",
INIT_09 => X"0820500B90419005B0C309402030060860E01004A828408800440405E3502940",
INIT_0A => X"A2020010100007865421432121804021C20452880C2D200000045C18C0E0000A",
INIT_0B => X"371097006026226495446E2110AE4417411204400000306B8186185C42900693",
INIT_0C => X"A00308003080030800308003080030800308001840018400400602A018809800",
INIT_0D => X"4008081010108003C000210020460801001FB3650C50DB13111C0D95C20C2030",
INIT_0E => X"14804032007E281F840C00284A17210001060D8306C18360C1380A0260CB9808",
INIT_0F => X"1555D5D79BBEF8E50B041029075982BF3873041029079982BF39748AA0AC8000",
INIT_10 => X"5156AEA479BFD7F7F3041029075982BF3E73041029079982BF3F632C5F96D3C1",
INIT_11 => X"932C5F96A595405FC7F1CFEBC7586C4100A53162B47FD7E39FFEECE159870234",
INIT_12 => X"39464006FE037ACFB88083A99E06271BB0CA207DFDD5920057E0B001B0EBCC79",
INIT_13 => X"6F5DF5CA2A002DD51B6F7FC4A411D1E8D44517F14EAFE36E55150016EA8DB73E",
INIT_14 => X"9DB84953C30351452A13D55CFFA76E928E3891F148B30399F5FB7F28C800DFA0",
INIT_15 => X"110155AC57DFEAEF1005475F1D1F608819CF0EE76E12C824ADD9089715F25FAF",
INIT_16 => X"0D8360D834041A41A0000010180C02801680460FC900052FA10DC0006DA4881C",
INIT_17 => X"D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D836",
INIT_18 => X"8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360",
INIT_19 => X"B000000000000000000000000020D8360D8360D8360D8360D8360D8360D8360D",
INIT_1A => X"1451451451448982C8A82E0820825942495377D9D701DC2E784601F8D187BEF8",
INIT_1B => X"4A2512A954AA5528944A25555145145145555555145145145555555145145145",
INIT_1C => X"FFC00000944A25128944A25128944A25128944A25128944A25128944A2512894",
INIT_1D => X"A5D2E820BA550000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFBFDFEFAAD142010007BEAB55FFAA821FFFFFFFFFFFFFFFFFFFFF7FBD74A",
INIT_1F => X"1FF002A821FFFFFFFFFEFF7D16AB55A2D542000A2D5400BA0800021FFFFFFFFF",
INIT_20 => X"DFFFFFFFC0010F7842AA10F780021FFFFFBFDF45A2D56AB45FFFFD54BAFF8000",
INIT_21 => X"6AB45A28000010082A975EFA2D140145007BC21FF5D2AAABFFF7D168B45AAD57",
INIT_22 => X"BC214555003DE10A2FBEAA00000002010552E95410AAFBD75FF5D7FEAB550051",
INIT_23 => X"04174AA5D00020BA555542145A284155FF5D517FE000004020AA552E80000F7F",
INIT_24 => X"00000000000017400082E954AA0800154AA0855575FFAAD57FE005D7BD740008",
INIT_25 => X"FFFFFDFEFF7FFD74AA552A820AA490A000000000000000000000000000000000",
INIT_26 => X"A080A051FFFFFFFFFEFF7F1FAFD7A2D5400001C7BEDB7DEBA4871FFFFFFFFFFF",
INIT_27 => X"6DFFFBD54AAE38E021FF0824821FFF7F1F8FC7EBD568B7DB6DF47000AADF400A",
INIT_28 => X"BC7E3D56AB7DB6DF78FD7EBF1C2000F78A2DA38E38A021C7E3F1F8F55AADB6FB",
INIT_29 => X"25EF497FEAB7D145B6FB45AA8E070281C20925FFBEDB451451C7BC01EF4124AD",
INIT_2A => X"00092412A87010E3F5C0145410E3DE28B6FFE8A101C0E05010412495428AAF1D",
INIT_2B => X"B7AE385D7FD74381400124825D0A000BA555F47145BE8A105EF555178E381C0A",
INIT_2C => X"00000000000000000000000000000154280024924AA1404174AA0055505EFBED",
INIT_2D => X"A80155FFFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA082A8000000000000000",
INIT_2E => X"F7FBD5410AAFBC00AA002A955FFF7FBFDFEFFFD568B45AAD5400005D7BFFFEFA",
INIT_2F => X"5AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF0000021EFF7D16AB55A2D56ABEF",
INIT_30 => X"45557BC21FF08003FF55AAD168BFFF7FFEAB45AAD140010F7AABFEBAAAAA8214",
INIT_31 => X"4100000154AAA2D1421FF007BE8BFF557BFDF55A2AA974AA5D04001EFFFFFD55",
INIT_32 => X"01EF55516AAAA5D2A82000082E95400A2D542155002ABDEBAF7FBE8A00552E95",
INIT_33 => X"174AA0855421FFFFFBEAAAA5D7BD74BA5D0002010552E820AA5D7BD7545F7AA8",
INIT_34 => X"0000000000000000000000000000000000000000000000174BA0004000AA5500",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000001000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000008128000000000000000000000024001620280000000000354200004008",
INIT_04 => X"000058800004C4024024001210001054B1C822009640000E2000002604003000",
INIT_05 => X"07008000E0200000000000000000200604000000001C04000026400000002C40",
INIT_06 => X"000000000000000004C010B35420015040000000002C42010010200004C83810",
INIT_07 => X"06E200201C00A14080082B26208008A009001201014022404402800408408020",
INIT_08 => X"00004180261C81210031000004340000200008105428020568040213003499C0",
INIT_09 => X"0000000990000000B0C308000000000860200160000000000038380000000000",
INIT_0A => X"10000000000005860000000080A0002060204080000000000004540800000000",
INIT_0B => X"00000000000000020001000022000000000000000000178000F8000101259000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000108000EC000000000000000010004B200000000000000000000000000",
INIT_0E => X"2000000000062801800400000000000000000000000000000000000000000000",
INIT_0F => X"828008084451B81A70AB3006BA0011400760AB3006BA0011400680F020968348",
INIT_10 => X"30B8011204082248A0AB3006BA0011400160AB3006BA0011400084C780687DBA",
INIT_11 => X"64C78068796E80A00802301BC0A7531EDD98E73B02800804620D030F873EB49F",
INIT_12 => X"B0A936B00000002044F091A860700FF9198AA115D5DA37F7A80C8A3604001C06",
INIT_13 => X"0000098551AC9000000000314E01F9F30198600631448410A2A8D64800000081",
INIT_14 => X"1046B2E00303842281C80A23004411AD661891F15148A4420804241526D60000",
INIT_15 => X"66A4A9D335F3D282000C6C5456C84850F61050C411AD6284FDA861682805A04A",
INIT_16 => X"0000000000000000000000000000000000004600C00138000030880042023043",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"9000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C30C30C30C3451046260A9A69A603924554117747E18E0218CC01400163A20C",
INIT_1B => X"26934984C26130984C26130C30C30C34D30C30C30C30C34D30C30C30C30C30C3",
INIT_1C => X"FFC000004C26130984C26130984C26130984C26130984C26130984C26130984C",
INIT_1D => X"A5D2A800105D2E80000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFF7FBD74AA5D2E820BA55003DFFFFFFFFFFFFFFFFFFFFFFFFFD54A",
INIT_1F => X"B55FFAABDFFFFFFFFFFFFFFFFFDFEFF7FFD54BA5D2EA8BFFFF84021FFFFFFFFF",
INIT_20 => X"8B55A2D540010007BEAABAA2AE821FFFFFFFFFFFFFFBFDFEFAAD142010007BEA",
INIT_21 => X"021FFFFFFFFFEFF7D16AB55A2D542000A2D5400BA08003DFFFFFFFFFFFFF7FBE",
INIT_22 => X"FD54BAFF80001FF002ABDFFFFFFFFDFEFA2D56AB45AAFBD74AAFFD5420100804",
INIT_23 => X"FBE8B45AAD568BFFF7FBD74BAFF802ABFFFFAE821FFFFFBFDF45A2D56AB45FFF",
INIT_24 => X"0000000000002ABFFF7D168B45AAD57DFFFFFFFC0010F7842AA10F780155FFF7",
INIT_25 => X"FFFFFFFFFFFFBD54AA5D2A80000412A800000000000000000000000000000000",
INIT_26 => X"7E384071FFFFFFFFFFFFFFFFDFEFF7FFD74AA552A820AA490A38FFFFFFFFFFFF",
INIT_27 => X"D7A2D5400001C7BEDB7DEBA4BAFFFFFFFFFFFFF7FBFDFD7EBF1D24AA5D2AADBD",
INIT_28 => X"FFFFFFBFDFC7E3F5EAB45AAD140000007FEFA92A2AA851FFFFFFFFFEFF7F1FAF",
INIT_29 => X"74AAE3DF400000004021FFF7F1F8FC7EBD568B7DB6DF47000AADF400AA080A3F",
INIT_2A => X"F8F55AADB6FB6DFFFBD54AAE38E021FF0824BDFEFE3F1F8FD7AAD16DB7DBEFBD",
INIT_2B => X"A2DA38E38A125C7E3F1EAB55B6DB6FBD7E3F5D04AAFF8A2DBD7E3A0821C7E3F1",
INIT_2C => X"000000000000000000000000000002DBC7E3D56AB7DB6DF78FD7EBF1C2000F78",
INIT_2D => X"82AA8BFFFFFFFFFFFFFFFFFFFFF7FBD54BA552A80010002A8000000000000000",
INIT_2E => X"A2D5400AA552ABDF55A280155FFFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA0",
INIT_2F => X"FF7FBFDFEFFFD568B45AAD5400005D7BFFFEFAA8028BFFFFFFFDFEFF7FFFFF55",
INIT_30 => X"10AAFBC00AA002ABDFEFF7FBFDF55AAD16AB55AAD140010007BFFE10AAAA955F",
INIT_31 => X"B45A2D57DFFFFFFFD54AAA2FBC20100800021EFF7D16AB55A2D56ABEFF7FBD54",
INIT_32 => X"FF45AA8002145AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF00003FFEFA2D56A",
INIT_33 => X"EAB45AAD140010F7AABFEBAAAAA82155AAD568B55FFFFFDF55A2D1400AAF7AAB",
INIT_34 => X"00000000000000000000000000000000000000000000003FF55AAD168BFFF7FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000002000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"000079800014CC02C034001600000000000000101EC0012EE0C0026E1E80F000",
INIT_05 => X"1F0FF433EFF0440C3902100002203F2EFC040388137C3E20C8EEC00284033CC0",
INIT_06 => X"7000660016490201700000000002FF57C8E8840155FDC0000010E40087D8787A",
INIT_07 => X"4000040007700000000000000001080FF900160000000200C00080001840BFE4",
INIT_08 => X"0009FFBFE5181606000410A4000004202AA8043E0000000000000001209244C0",
INIT_09 => X"0001227FB0000000F7DF78020004011FEFE00000000020031502000083880200",
INIT_0A => X"00000000000015BE0000004000000100000100506002008C2007D5FC80000024",
INIT_0B => X"0020000000000000000000000000000000210018800000000000000010000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000020",
INIT_0D => X"0008000000100000010000002000080101FFB600000000000000000000000000",
INIT_0E => X"0000003007FE29FF800C00000001002040000000000000020480002E42429C00",
INIT_0F => X"000000004D4E180010040000400000001E60040000400000001E6010003C0000",
INIT_10 => X"04000000000094B1E0040000400000001E60040000400000001E608040000004",
INIT_11 => X"0080400002000000000033628000100100000004000000006170C00080010000",
INIT_12 => X"B0020000000000295810000000A100020614148002000000000004307CC3CC00",
INIT_13 => X"000525802000000000014AC000120200000000003F0D800020100000000000A4",
INIT_14 => X"000020020C0C00000000002E2D000001006204040000000005786C0040000000",
INIT_15 => X"004000100A0C0939BEE1810080200000E0CE0EC000010020000000000000AE8A",
INIT_16 => X"000002008040400400C08080000000000049F6FFC01000000000000080080080",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"6902001000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"186186186190324C1090D0F3CF3CD039A060000600704000201120AB02090082",
INIT_1B => X"0C86432190C86432190C86596596596596596596596596596596596596596186",
INIT_1C => X"FFC00002190C86432190C86432190C86432190C86432190C86432190C8643219",
INIT_1D => X"A552A82010080400000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD54AA5D2A800105D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"0BA5500001FFFFFFFFFFFFFFFFFFFFFFFBD54BA552A8001000003DFFFFFFFFFF",
INIT_20 => X"FFEFF7FFD74BA552E801FF002E821FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E82",
INIT_21 => X"BDFFFFFFFFFFFFFFFFFDFEFF7FFD54BA5D2EA8BFFFF843FFFFFFFFFFFFFFFFFF",
INIT_22 => X"142010007BEAB55FFAA801FFFFFFFFFFFFFFBFDFEFFFD542000082EAAB55AAAA",
INIT_23 => X"FFFFFFFF7FBFDF55AAD140000087BE8B55F784021FFFFFFFFFFFFFFBFDFEFAAD",
INIT_24 => X"0000000000003DFFFFFFFFFFFFF7FBE8B55A2D540010007BEAABAA2AE975FFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA552A820001400000000000000000000000000000000000",
INIT_26 => X"81C0038FFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2A80000412ABFFFFFFFFFFFFF",
INIT_27 => X"EFF7FFD74AA552A820AA490A021FFFFFFFFFFFFFFFFFFEFF7FBD74BA5D2A8002",
INIT_28 => X"FFFFFFFFFFFFFFFBFDFEFFFFFD54BA5D2A801C7142E871FFFFFFFFFFFFFFFFDF",
INIT_29 => X"0010142AAFB7DBEAEBAFFFFFFFFFFFFF7FBFDFD7EBF1D24AA5D2AADBD7E38438",
INIT_2A => X"FFFEFF7F1FAFD7A2D5400001C7BEDB7DEBA4871FFFFFFFFFEFF7FBF8FD7E3D14",
INIT_2B => X"FEFA92A2AA925FFFFFFFDFEFE3F1FAF45A2D142010087FEDB55F78A051FFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFBFDFC7E3F5EAB45AAD140000007",
INIT_2D => X"02ABFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005D040000000000000000",
INIT_2E => X"F7FFD74AA5D2A800BA550428BFFFFFFFFFFFFFFFFFFFFF7FBD54BA552A800100",
INIT_2F => X"FFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA082A821FFFFFFFFFFFFFFBFDFEF",
INIT_30 => X"AA552ABDF55A2802ABFFFFFFFFFEFF7FBFFFFFF7FBD74BA552A80145552E955F",
INIT_31 => X"FEFF7FFEAB45AAD1420105D2ABFFFFFFAEA8BFFFFFFFDFEFF7FFFFF55A2D5400",
INIT_32 => X"DF55F7AE955FFF7FBFDFEFFFD568B45AAD5400005D7BFFFEFAA80175FFFFFBFD",
INIT_33 => X"6AB55AAD140010007BFFE10AAAA821EFF7FBFDFFFAAD168B55A2D542010007BF",
INIT_34 => X"00000000000000000000000000000000000000000000003DFEFF7FBFDF55AAD1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"084A76341244919000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"000079800014CC03C075161E001118653D2408041FC004AEF000816E1C11F541",
INIT_05 => X"3F0F807BFFE000240100004683103E7FFE02482553FC3C0204EFC25010143CC0",
INIT_06 => X"1100441004201014B1709C910102FF5FC0A0000101FFE4036450E08247F87870",
INIT_07 => X"08750504800680102542AD800504530FF9061E8026998E9A00402CC25BD0FFFC",
INIT_08 => X"0011FBFFE04691A5A00101818A6800088228000001A044C8168480D010F200AA",
INIT_09 => X"B6E85A7FF080AC70FFDF78220010841EFFE7116E144071268DFD3E4C24040100",
INIT_0A => X"3151518A8A31B7FE00040009814C089202225412115428C03BC7D7FC15025B1A",
INIT_0B => X"1B1883007104032901CC63410ABD249C4B338934404037FC8BFE18008083B444",
INIT_0C => X"D9228D9228D9228D9228D9228D9228D9228D99146C9146C84006309044081A00",
INIT_0D => X"48000201800500941044312000900D4621FFBE00080081529904595123203040",
INIT_0E => X"308162029FFEADFF8050250010030165290008800440022201082401A002000C",
INIT_0F => X"5001318048A004A6C0D2820302C005A83480D1820302A009B02B101390C0CB28",
INIT_10 => X"485101408904831400D1820302C005A83480D2820302A009B02B021A85C09411",
INIT_11 => X"FA1A85C08834600024D052C1051E0B92D400360520202682C19024B6164E3004",
INIT_12 => X"C1B0D6404093E22A2012418A9D1D44ADD9E0F174103820101C0B8160D5516259",
INIT_13 => X"6C88660D8AA288209E615100280DA0052000C5006402000206C55144104D510C",
INIT_14 => X"024500A0D50020C04023033C52009144231D902818100C90058010361AC80812",
INIT_15 => X"198A12202386454988140600C0181500A13E830011008B0374007000B4E0CD00",
INIT_16 => X"008020080224004002000000703804008001F7FFF01B982B01258088C008CC41",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"F000000000000000000000000020080200802008020080200802008020080200",
INIT_1A => X"7DF7DF7DF7DFFFFEFEFFFE79E79FFFF3BC1FF3FDDFEFFFBEFFE7DF84081EFEFB",
INIT_1B => X"FEFF7FBFDFEFF7FBFDFEFF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF",
INIT_1C => X"FFC00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"A5D2E80010000400000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA552A8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"0105D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E80010552EBFFFFFFFFFFF",
INIT_20 => X"FFFFFFFBD54BA5D2E82010002ABDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A80",
INIT_21 => X"001FFFFFFFFFFFFFFFFFFFFFFFBD54BA552A800100000001FFFFFFFFFFFFFFFF",
INIT_22 => X"BD74AA5D2E820BA5500001FFFFFFFFFFFFFFFFFFFFF7FBD74BA5D2E800BA5D00",
INIT_23 => X"FFFFFFFFFFFFFFEFF7FBD74AA552A800BA5D2E821FFFFFFFFFFFFFFFFFFFFF7F",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFEFF7FFD74BA552E801FF002E975FFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E800000800000000000000000000000000000000000",
INIT_26 => X"05D2ABFFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8200014003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFBD54AA5D2A80000412ABDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2E8000",
INIT_28 => X"1FFFFFFFFFFFFFFFFFFFFF7FBD54BA552E82028002AB8FFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74AA5D2E800AA5500021FFFFFFFFFFFFFFFFFFEFF7FBD74BA5D2A800281C0000",
INIT_2A => X"FFFFFFFFFFDFEFF7FFD74AA552A820AA490A071FFFFFFFFFFFFFFFFFFEFF7FBD",
INIT_2B => X"A801C7142E955FFFFFFFFFFFFFFFFDFEFF7FFD54BA5D2E80082492E871FFFFFF",
INIT_2C => X"0000000000000000000000000000038FFFFFFFFFFFFFFFBFDFEFFFFFD54BA5D2",
INIT_2D => X"D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008000000000000000000",
INIT_2E => X"FFFBD54AA5D2E800005D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF7FBD54BA552A80010002ABDFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"AA5D2A800BA5504021FFFFFFFFFFFFFFFFDFEFF7FBD74AA552E820BA002AA8BF",
INIT_31 => X"FFFFFFBFDFEFFFFFD54BA552E800BA5D04021FFFFFFFFFFFFFFBFDFEFF7FFD74",
INIT_32 => X"0000082A955FFFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA082A955FFFFFFFF",
INIT_33 => X"FFFFFF7FBD74BA552A80145552E975FFFFFFFFFEFF7FBFDFFFFFFBD74AA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000002ABFFFFFFFFFEFF7FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"431965109E4481D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"492C0020220001010E4916C884DCD607E5EC2A344103E48003D0800023D0072C",
INIT_05 => X"00107C441001100D620A06D683018001023D37E5088043620101179092540112",
INIT_06 => X"401002010042384D223C19C3552800081ADA0E054402365774611E047020008E",
INIT_07 => X"491EC04ED017AB5497EB923F08182E20020689B735011FBFE7BC062602944019",
INIT_08 => X"154A00401D4425ADA9035BE19C8F9442A8801200F4C9D7AC8093A051727B2AC3",
INIT_09 => X"9A50020040E48D50080002B00A0C00801014541E9504703680017F6CB4050700",
INIT_0A => X"8151538A8A738041C23020131A80CFDFF3FE509A907C6AC05040220409009031",
INIT_0B => X"2D040050110081E9528963546278008AA80381B4000500026800000109379864",
INIT_0C => X"1C2A81C2A81C2A81C2A81C2A81C2A81C2A81C9540E1540E00140000610000320",
INIT_0D => X"594A06870A9CA0D458D131652A154D46B6000850800801628013456520CA0928",
INIT_0E => X"02080448C00044000A1EC1C44140D101A54280A14050A028500A84F02842A24C",
INIT_0F => X"0061338359E0C4E6C256690581800F1C3E82562B0581200F1C3F081456022804",
INIT_10 => X"2C438100AB8581B602562B0581800F1C3E8256690581200F1C3F1238473F1210",
INIT_11 => X"2238473F0E1050083750B3E4275F829547008600C030374361FA2CEE046D4812",
INIT_12 => X"C1128C4CC012A66F61154C019511628756231018500C00203E13806156516078",
INIT_13 => X"54CDE608AA612C0096C37B00D1724801A0009C606D1221D104553096004B61BC",
INIT_14 => X"870B012A41E0F0600035842E7601C2C4AC68A98810080AA825A8902251899802",
INIT_15 => X"58234A89637E00D0A1080301401C390320188321C2C0B13890105800D520AF94",
INIT_16 => X"8822088222F110111B281A54753AA004002601001918008C10912A4440B24E8B",
INIT_17 => X"8220882208822088220882208822088220882208822088220882208822088220",
INIT_18 => X"2008020080200802008020080200802008020080200802008022088220882208",
INIT_19 => X"E82891448000000001FFFFFFFFC8020080200802008020080200802008020080",
INIT_1A => X"3CF3CF3CF3DFFBFEFEBEEEFBEFBEFBEBFDF7F7FBDFD1FE3EFBD7ADFBF7EFBEFB",
INIT_1B => X"FE7F3F9FCFE7F3F9FCFE7F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"FFC00001FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"A5D2E82000000000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8000008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74AA552E8000055003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A82",
INIT_21 => X"BFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E80010552EBFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD54AA5D2A800105D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A82000552A",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD54AA5D2A800005D2EBDFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000000001FFFFFFFFFFFFFFFFFFFFFFFBD54BA5D2E82010002AA8BFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100004000000000000000000000000000000000",
INIT_26 => X"008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA552A8200014003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E800105D043FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"54AA5D2A82010552EBDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2E800005D2ABF",
INIT_2A => X"FFFFFFFFFFFFFFFFFBD54AA5D2A80000412AB8FFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E82028002AA8BFFFFFFFFFFFFFFFFFFFFFFFBD54BA552E80038492EB8FFFFFFF",
INIT_2C => X"00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFF7FBD54BA552",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000040000000000000000",
INIT_2E => X"FFFFD74BA552A8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E800000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005D043FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"AA5D2E800005D2EBDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA552E8001055003FFF",
INIT_31 => X"FFFFFFFFFFFFF7FBD54BA5D2A820105D2ABDFFFFFFFFFFFFFFFFFFFFFFFFBD54",
INIT_32 => X"00AA082EA8BFFFFFFFFFFFFFFFFFFFFF7FBD54BA552A80010002AA8BFFFFFFFF",
INIT_33 => X"FDFEFF7FBD74AA552E820BA002AAABFFFFFFFFFFFFFFFFFFEFF7FBD74BA552E8",
INIT_34 => X"0000000000000000000000000000000000000000000000021FFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"2C4360101A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"00017B810015DC03D034201E14000036486008101FC0002EE006297E1C05F561",
INIT_05 => X"BF0F817FFFE80100004044800080BEFFFC0248005FFC3C18A5FFC2444484BCC0",
INIT_06 => X"B0801408110000109127E0500002FFDFC000000001FFC0832050E00047F97870",
INIT_07 => X"00D1D72040048D00388387D03D0E591FFD201F862691DFBE077C2BC45B40FFE4",
INIT_08 => X"001FFBFFEC440501A5604B31062356282AA84200D12342113EDC400000045828",
INIT_09 => X"25A890FFF0002023FFDF79000000000EFFE309606020008005FC000000402000",
INIT_0A => X"30000000000037FF50010103134CAFDF03BA18000F39A0106F87D7FA84024B02",
INIT_0B => X"1B188300624483890564084198AD249C43300C00415037FC83FE1840C0902400",
INIT_0C => X"C1010C1010C1010C1010C1010C1010C1010C10086080860840063090442A1800",
INIT_0D => X"0001403000100200180480000095280001FFBF040C40C81119A41C1443243050",
INIT_0E => X"32A163821FFEAFFF805025E00853B92588000400020001000020A80180080020",
INIT_0F => X"90401486148484054395E27E428002A4200397E07E422002A420100382FCC308",
INIT_10 => X"641100C0788417000397E07E428002A4200395E27E422002A420110A51C01C05",
INIT_11 => X"C90A51C01A2490040590C08120558C1759BE1C05A0400383808800DA1929F728",
INIT_12 => X"00CE720000136006000215EA0A4833A32C8832050028603050014031B3950000",
INIT_13 => X"6C00C006658280009A2030108B14AC05C00112405222088B8332C140004D1018",
INIT_14 => X"A2659196B6808060201281004228996085F10020180C030880D11019CE400002",
INIT_15 => X"0108152A49DC7143F01C04240030720641E0A028996483A17204680410A04104",
INIT_16 => X"040100401000080080000000000002001201F7FFC0011C2F81A48080CA32800A",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_19 => X"0000000000000000000000000000401004010040100401004010040100401004",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000020000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFC0000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2A8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E80",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8000008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA552A8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A820000004",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA552A8201000043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E8000055003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA552A8200008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001008043F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA552A8200014003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E800105D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E820101C003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552",
INIT_2D => X"0043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA552A8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001008043FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74AA552A8200008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"200055043FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005D043FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD54AA552E8001055003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA552E8",
INIT_34 => X"00000000000000000000000000000000000000000000003DFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"00003A2E200811000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"000079800014CC03C034001E04010850300000101FC0002EE000006E1C00F500",
INIT_05 => X"1F0F8033FFE000000000000000003E2FFC024800137C3C0000EFC00000003CC0",
INIT_06 => X"000000000000000091C115500002FF5FC000000001FFC0000010E00007F87870",
INIT_07 => X"10E600084002040A10812A000500590FF9001F95406A8000037230C01840FFE0",
INIT_08 => X"0001FBFFEC4695A501604A000C7585080002C200408102F16C0184800026C92C",
INIT_09 => X"24A8107FF0000000FFDF78000000000EFFE001600000000005FC000000000000",
INIT_0A => X"30000000000037FF4000000AA0354000019C4000012800002387D7F804024B02",
INIT_0B => X"1218830060040A04000400000801241443300800404037E883FE180000000000",
INIT_0C => X"C1000C1000C1000C1000C1000C1000C1000C1000608006084006301044081800",
INIT_0D => X"00000004800B0000000000000000000001FFBE00080080101904181003003000",
INIT_0E => X"B08062021FFEADFF800020800000002088000000000000000000200180000000",
INIT_0F => X"D0210840009181008024A00043601100210024A00043C0110020901382CCCB28",
INIT_10 => X"0C920180040A03080024A00043601100210024A00043C01100209240C840C201",
INIT_11 => X"1A40C840A604E0080820009908008341B000A821207008200289001006832086",
INIT_12 => X"0166B40600800082041205EC00044C1ACB66C37542082030281E058000101281",
INIT_13 => X"0010480B27A004300004103160DB3005E000618040C022000593D00218000209",
INIT_14 => X"880012BBFF20406040084210C062000C2A2DDD00180C04504086002CD680C010",
INIT_15 => X"4106020804295C98F80400008040CC0582169022000C2876C404780028500160",
INIT_16 => X"000000000000000000000000000000000001F7FFC001B823018F008800088052",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"C800000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"7CF7CF7CF7D933CC3090CABAEBAFF969319815DD5EDCF9822659AE7B095A220C",
INIT_1B => X"1E0F0783C1E0F0783C1E0F7DF7DF7DF3CF3CF3CF3CF3CF7DF7DF7DF7DF7DF7CF",
INIT_1C => X"FFC000003C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C",
INIT_1D => X"A5D2E82010080400000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"00000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E800000800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8001000003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100804000000000000000000000000000000000",
INIT_26 => X"000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"A8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000043FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008040000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8000008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"000008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2A8001008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00002000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"924279824C94CC1BE0B4001F20000000020380401FE0082EF000106E1C00F500",
INIT_05 => X"1F0F8033FFF048202582800100523E2FFE024820137C3C0040EFE02000003CE4",
INIT_06 => X"F10466105670019C900000100002FF5FC0E0801101FFC0000010E08A07FC7870",
INIT_07 => X"0000040000000000000000000500590FF9001F0000000000033020C01840FFFC",
INIT_08 => X"0001FBFFFD0004000100502000011400000282004001020000000001009015C0",
INIT_09 => X"2CB8DA7FF8004000FFDF7C062031863EFFF75D78004001010DFC000020050100",
INIT_0A => X"30000000000037FFC00602000000000001980400002800032387D7FE94FBEF2B",
INIT_0B => X"9258830060040200000400000801243443B00808404037E883FE180C00000000",
INIT_0C => X"C1000C1000C1000C1000C1000C1000C1000C10006080060840077330C4889CC2",
INIT_0D => X"0000000000000000000000000001280001FFBE00080080101904189003003000",
INIT_0E => X"30A063021FFEADFF805025C0304001E58906088304418222C108A009A0904000",
INIT_0F => X"1000000000100100000480000200100000000480000200100000100380F0C308",
INIT_10 => X"0010000000080000000480000200100000000480000200100000000040400000",
INIT_11 => X"0000404000040000000000080800000110000000200000000200000000012000",
INIT_12 => X"00021000000000800002018C0100000208000008001220000000040040000080",
INIT_13 => X"0010000020800000000400000010200200000000008002000010400000000200",
INIT_14 => X"0800000210000080010000008002000000210000201000000002000042000000",
INIT_15 => X"0184000000084000000006050000000002000002000000204000000000000020",
INIT_16 => X"08822288226410410346010000000400A011F7FFE00318230104008000008000",
INIT_17 => X"8822088220882208822088220882208822088220882208822088220882208822",
INIT_18 => X"8220882208822088220882208822088220882208822088220882208822088220",
INIT_19 => X"0404000017FFFFFFFFFFFFFFFFE0882208822088220882208822088220882208",
INIT_1A => X"492082492085048029890AD34D35FDD04A165129432D518B45265EFC30760AED",
INIT_1B => X"C46231188C46231188C462492492492492492492492492082082082082082082",
INIT_1C => X"FFC000058AC562B158AC562B158AC562B158AC562B158AC562B158AC562B158A",
INIT_1D => X"A5D2E820100800000000000000000000000000000000000000000000000003FF",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100000",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000043FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"4A53D958C50000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"DBFAFBD7FB1CDEBEF1BE17F7AC88042787FBFFF8FEE9FF7EE6F4C0EE1FFAF869",
INIT_05 => X"5F0FFEB3EFFEFFBDA7F7FED508707E2EFEBF6FFEB37C3FF302EEEDFF9B487CF6",
INIT_06 => X"74EADE4EBDFDAC9930F6F8129E3FFFF7C3E3A74667FDDB7FB870FF30FFDEF87F",
INIT_07 => X"8173840C07783060C72DF7D828912E6FFB80162776F3BFB7077E82255E40BFEF",
INIT_08 => X"4769FFBFE43C872321367036163F1C0820A3063F460D1AEFC000060042648C41",
INIT_09 => X"BEFB967FBD13D981F7DF7D7E6171AF3FEFE8A3E679FAC1FD1FFFBEB000763A84",
INIT_0A => X"F3A3AD1D1DAD7FBE7D67D7F3BB79CFFB83BF14EC1E7D7300B017F5FFE6FBEF73",
INIT_0B => X"52199F58F6EE6F5E7FAC4C03DB856CD4CF720FE8C4427FF8CFFE38FF7F6BD928",
INIT_0C => X"F78C0D78C0D78C0D78C0D78C0D78C0D78C0D7A606BC606B8C56F7730ECCDBDF1",
INIT_0D => X"EA035CF6100C0E60FB9FC3A80EF69A04DFFFF7FF5E75FF341B867D3683A03A40",
INIT_0E => X"36B867027FFFF9FF8FAFAA3ADEBFB9726BAF5FD7AFEBD7F7EFFD7ACDB7F947F0",
INIT_0F => X"10003E020080A40403E8BD8002000FC02003E8BD8002000FC02010979AFFE36C",
INIT_10 => X"80100000EE00034003E8BD8002000FC02003E8BD8002000FC020037B0040A000",
INIT_11 => X"037B0040C00400003D80008160400FD81341C00020003B80008C00801EF02853",
INIT_12 => X"01F1190981038406809677FA080468C46A81080581002000780C8001C8100201",
INIT_13 => X"7080D00F90D162001C803411FC0024080001F80040026C0807C868B1000E401A",
INIT_14 => X"B02013F810503A00003E020042AC080CEB01228A80000F600080123E23213040",
INIT_15 => X"61F810087520750001064180807868000110C02C080CFA0042400000F8800105",
INIT_16 => X"5FD7F7FDFF7EFEEFF3EEC3FF7FBFFBCB7FFFFEFFE00BFF7FEBF420800EC0CBEE",
INIT_17 => X"FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F",
INIT_18 => X"D7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5",
INIT_19 => X"6DAE443237FFFFFFFFFFFFFFFFF5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5F",
INIT_1A => X"4D34D30C30DD795EAA6AFC38E38EA3AB788962B79E923C2CD990A7D3B4A9FC37",
INIT_1B => X"26130984C26130984C26130C30C30C30C30C30C30C30C30C30C30C30C30C30C3",
INIT_1C => X"FFC000004C26130984C26130984C26130984C26130984C26130984C26130984C",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"0842D85841000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"DBEAE5D6D91C2EBCE1B21EA72C00000007FBE7C8F8E9EF79E6D440E91FDAE061",
INIT_05 => X"5C8FFCB38FF6B68984B5BCE408347E28FEBF6FEEB3723F7102E8EDBF8A4872F6",
INIT_06 => X"946ACF46ACE0841A00006A089E3FFF27C3032646EFF1DB7FA868FE30EF1CE47E",
INIT_07 => X"8000000A20083060C00C81882A008C6FF880060424B39FB6037F00051C003FE0",
INIT_08 => X"4761FA3FE4010440410844060001040A00002200460D1A060000050400000010",
INIT_09 => X"FEEB027E390A4881C7BEFC5F6171CE2F8FE823E778DAC16C1FFBBC9000315895",
INIT_0A => X"F606013030213C3E2D62D6E21259CFDB039E806C024531008017C1F826FFEF41",
INIT_0B => X"5219AB5AF86F7D5E382A440349816DD4C7560B60D4427FF0C7FEBABF3F6BD108",
INIT_0C => X"E3440C3440C3440C3440C3440C3440C3440C3C2061A2061AD46FF730E5CCBCD5",
INIT_0D => X"6203E8FC10080A20ED1D41880CC61A044DFFC6EB5AB5B7941BC63F1683803C00",
INIT_0E => X"B88572023FFE91FF98AEAA1AC6AC9A3A4AAD5B56ADAB56D5AFD572C597B14750",
INIT_0F => X"10003E020000260403C8948002000EC0000BC8948002000EC00010878AC3CB8A",
INIT_10 => X"80100000EE0000400BC8948002000EC0000BC8948002000EC000097B00402000",
INIT_11 => X"017B0040400400003D80000070400DD81041400020003B80000410801AF02041",
INIT_12 => X"05D11101010384008086378A080428C46A80080081002000780C800188000301",
INIT_13 => X"7080102E909042001C800409FC0020080001F80000007C0807484821000E4002",
INIT_14 => X"F02003F810100A00003E020000BC0808EB01020280000F60000002BA22202040",
INIT_15 => X"21F810007520750000024080807868000100403C0808FA0040400000F8800001",
INIT_16 => X"5B56D5B5EF3AF6AF6389C2FE128971AB2DDDF8FFE0031B776BF4208006C0C926",
INIT_17 => X"B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D",
INIT_18 => X"56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5",
INIT_19 => X"238B443A3FFFFFFFFFFFFFFFFFD5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B",
INIT_1A => X"00000000000F0080397908000000A4805F09C42D0200903950C086D420010825",
INIT_1B => X"8040201008040201008040000000000000000000000000000000000000000410",
INIT_1C => X"FFC00005028140A05028140A05028140A05028140A05028140A05028140A0502",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100804",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"461080404900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"00800040110102000902002000888400081045A8A00003C00000500000080008",
INIT_05 => X"0000000000024CA0A0101800032000400000000B800000014000000B08180000",
INIT_06 => X"0020280202802C00020800008A14002011110012220009A88800009A88000000",
INIT_07 => X"8108044200091224484510201000204000800020410000000080000104000009",
INIT_08 => X"132800000140200808021006108010422AAA8000224489028492201140092240",
INIT_09 => X"0001C800004080A0000002480B04008100011000088800081002C19020150B00",
INIT_0A => X"4353529A9A528000040040702080000000400064080011001050000200000018",
INIT_0B => X"01400048012220122A0004168110400004000040811600000400001036584108",
INIT_0C => X"36050160501605016050160501605016050160280B0280B00120008430660210",
INIT_0D => X"2A000C4210040860B188C0A8065302005A0040390010120500002002C0040010",
INIT_0E => X"8221050060001000028000080205001066000100008000400490020402010530",
INIT_0F => X"000000000000A00000081480000001400000081480000001400000800C010820",
INIT_10 => X"8000000000000240000814800000014000000814800000014000000100002000",
INIT_11 => X"000100004000000000000001400000080041400000000000000C000000100041",
INIT_12 => X"000101010100000480802A400000004000000800810000000000000048000000",
INIT_13 => X"0000900010104200000024000400000800000000000244000008082100000012",
INIT_14 => X"1000004000100A00000000000284000040000202800000000000120020202040",
INIT_15 => X"2050000010000000000240800000000000104004000040000040000000000005",
INIT_16 => X"010040108408420430E699AA42A1508104EA08000000810020000000044001AC",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"0506117080000000000000000000100401004010040100401004010040100401",
INIT_1A => X"4104104104006C1A8283AC618618EF10C0422205822140048D2E581E80DEC4D2",
INIT_1B => X"C06030180C06030180C060410410410410410410410410410410410410410410",
INIT_1C => X"FFC0000582C160B0582C160B0582C160B0582C160B0582C160B0582C160B0582",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0401D940CD0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"49B87A417315D20A313E17F1800000058013DDF8BE21F36E02F0D06E03E8F800",
INIT_05 => X"1F007E33E01A4D9C87525E5101603E6E023D27DA937C03E340EE25CB9B483C12",
INIT_06 => X"F0A05A0A15AD0C0130F6F0128A16FFF001E1870223FC3BFC98101F109FC6780F",
INIT_07 => X"8073800407781020476467D008910A4FFB80100332D1AE93059282215E408006",
INIT_08 => X"0221FF80003C832320342036063F08000001063F42050AEB4000221000248C01",
INIT_09 => X"9A51547F8C1111A0F041056A0100A11FE000916249A800B915FE82B020522900",
INIT_0A => X"42A2AD1515AD5780540541619968C76980E914E4163D53002017F405C409A42A",
INIT_0B => X"0140140816A22B126DA40C03531440800C2005C8800217F80C000055FF7C4928",
INIT_0C => X"268D0068D0068D0068D0068D0068D0068D006A68034680300021410028450530",
INIT_0D => X"AA01587410080C60AB0F42A804628200DBFFF13D04505B2500806522C0A40A50",
INIT_0E => X"941922006FFFF8000F8F80281A16A1504302058102C0816244B82A0CA25907D0",
INIT_0F => X"000000000080A40000283D80000001402000283D80000001402010901A7D6944",
INIT_10 => X"800000000000034000283D80000001402000283D80000001402002010000A000",
INIT_11 => X"02010000C000000000000081600002080341C00000000000008C000004100853",
INIT_12 => X"0021090981000006809076B20000404000010805810000000000000048100200",
INIT_13 => X"0000D0011051620000003410040004080000000040026C00008828B10000001A",
INIT_14 => X"B000104000503A000000000042AC00044000228A800000000080120421213040",
INIT_15 => X"607800081000000001064180000000000010C02C000440000240000000000105",
INIT_16 => X"05816258964C4A44A0C689FF3F9FFEC5D6DBFE0020096528A0B000000CC043EC",
INIT_17 => X"5816058160581605816058160581605816058160581605816058160581605816",
INIT_18 => X"8160581605816058160581605816058160581605816058160581605816058160",
INIT_19 => X"F506003017FFFFFFFFFFFFFFFFE0581605816058160581605816058160581605",
INIT_1A => X"5D75D75D75DFFFFEFCFDF7FFFFFF5DE7FC3DF3F2DDCFFFBEFFCF1F84421FFEFF",
INIT_1B => X"EFF7FBFDFEFF7FBFDFEFF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF75D7",
INIT_1C => X"FFC00007DFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDF",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"E800000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"3CF3CF3CF3DD7FDEBAFAFEFBEFBFFBFBB9DFF7FFDFF3FC3EFFF7FDFBBDFFFEFF",
INIT_1B => X"FE7F3F9FCFE7F3F9FCFE7F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"FFC00001FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"08425818000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"DB6A618248140C18E0B016872400000007EBA24058E1ECA8E2D400681FD0E061",
INIT_05 => X"1C0FFC338FF01009048084C400103E28FE3F6FE513703F7000E8E5B4825030F6",
INIT_06 => X"100046000460001800006800142AFF07C202060445F1F2572060FE82671C607E",
INIT_07 => X"00000008800020408008818838000C2FF800060424B39FB6037E000418003FE0",
INIT_08 => X"0441FA3FE4000400010040000001040880000200440912040000040000000000",
INIT_09 => X"BEE8027E38004801C79E7C162231862E8FE00166704041240DF93D0000000000",
INIT_0A => X"B00000000000343E002202021259CFDB039E0008024520000047C1F804FBEF01",
INIT_0B => X"121883107044094C1028400548812494C3120920404437F0C3FE180D89279000",
INIT_0C => X"C1000C1000C1000C1000C1000C1000C1000C18006080060840477330C4889CC0",
INIT_0D => X"400340B400080200481501000884080405FF86400800811019861D1403803800",
INIT_0E => X"308062021FFE81FF880EA000400098200C04080204010200810020C180904240",
INIT_0F => X"10003E020000040403C0800002000E800003C0800002000E8000100780C2C308",
INIT_10 => X"00100000EE00000003C0800002000E800003C0800002000E8000017A00400000",
INIT_11 => X"017A0040000400003D80000020400DD01000000020003B80000000801AE02000",
INIT_12 => X"01D01000000384000006118A080428846A80000000002000780C800180000201",
INIT_13 => X"7080000E808000001C800001F80020000001F8000000280807404000000E4000",
INIT_14 => X"A02003B810000000003E020000280808AB01000000000F600000003A02000000",
INIT_15 => X"01A81000652075000000000080786800010000280808BA0040000000F8800000",
INIT_16 => X"08020080223010010308025410082404A015F0FFE003182701B420800280C802",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_18 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_19 => X"0008004017FFFFFFFFFFFFFFFFC0802008020080200802008020080200802008",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFC0000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"441406267B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"0005802424830120024121209088809DF81454ACA01E03501D0A3B91E00F0A00",
INIT_05 => X"E0F001CC00012034C20B0232838F80D001C0100AEC83C008EF101A034C8CC300",
INIT_06 => X"2F1620F1721BA346AA2C95C5CB1400000161F84322000DA8C40F003C80030780",
INIT_07 => X"5939F36677EE1C387777622717EF711004A6818111086008E080FDC305940018",
INIT_08 => X"13160400195E83A3A0F61BC3929ECB622AABF5FF83860CEB164833F179B48CEE",
INIT_09 => X"01036D8004FDB47600000229410C61010016DC998C84B0128202C0DCB48F05D5",
INIT_0A => X"4400402A0A37000182502440888420247041E876810099D35F900002DB00105C",
INIT_0B => X"AD4434020CA2E0B32B01A752B078412A24818094151348062400E2A034D86444",
INIT_0C => X"3E2781EA781E2781EA781E2781EA781E2781C33C0613C0E21028840239452116",
INIT_0D => X"394818429A95E954868AD0E52273F54258000080808900C3807122C3E04E0338",
INIT_0E => X"8E3B15C94001120055704DC4A1624487E2489024481224091282C4300942A194",
INIT_0F => X"C06101C55D65C3E3F01F52FFC1E0013C1F801F52FFC1E0013C1F8090423D38A1",
INIT_10 => X"ECC381C0118796BE001F567FC1E0013C1F801F567FC1E0013C1F9085DFBF7E15",
INIT_11 => X"F885DFBF7E30F00C0270F3751F1FD00FECBF7E25C0700463E17B2C7F811FD7AD",
INIT_12 => X"C40FE6474190626D6491063597F9177B956EF378D33E4030061341F077C571F8",
INIT_13 => X"0C4DAE207F328E3082636B2807FFD80FE00007E03F7207D3E03F9167184131B5",
INIT_14 => X"1F4FE047EFA0CAE06101C53E3647D3F144FCDD22B81C0098E57D9081FCE8C852",
INIT_15 => X"38574FF31ADF08DBF81846A540049707E0FE3307D3F141FFB45478040570EED4",
INIT_16 => X"90240902C189601208A1102B4AA5584B4068000019A80098120BCA4C617635C9",
INIT_17 => X"0240902409024090240902409024090240902409024090240902409024090240",
INIT_18 => X"2409024090240902409024090240902409024090240902409024090240902409",
INIT_19 => X"9AA09426A8000000000000000009024090240902409024090240902409024090",
INIT_1A => X"104104104104431042720EE38E38AAF9A93E7131C136AD8E9B562CF03B2E8E78",
INIT_1B => X"F87C3E1F0F87C3E1F0F87C104104104104104104104104104104104104104104",
INIT_1C => X"FFC00001F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0",
INIT_1D => X"AAAAABDEBAF7AE8000000000000000000000000000000000000000000000C200",
INIT_1E => X"EFF7D142145A2AE800BA08514214555517DEAA5D7BFFEAAF7803FEBAF7FFD74B",
INIT_1F => X"E00A2FBD75FFFF84001550851555FF55517FE000055421FF00557DF45A2D5401",
INIT_20 => X"74BA552EBDFFF0004020005D5555555A2AABFFFF5D516AA00A28028A00AAAEBF",
INIT_21 => X"3FEBA082ABFE10AAAEA8ABA55517FF45A2AEBDEBAAAAAA8BFFF7D140010FF841",
INIT_22 => X"FD75FF0051401FF5D00154105504000BA5D2E97545A28028B450855401450804",
INIT_23 => X"FBFFF45A2FFFDE00002E801FFA2AABFE00FFFFD74AA085540000002E801FF557",
INIT_24 => X"0000000000002ABEFAA80001EFF7FFC20BAF7D1575450800020BA08517FF45F7",
INIT_25 => X"57803AEBAF7F5D74AAA2A03AA38BF8FC00000000000000000000000000000000",
INIT_26 => X"7A3F00516DA2D5451D7EBDB47155BC2A87092AAFA9257F1C5BC00AA5D7FF8EAA",
INIT_27 => X"00EA8000150A801C01C7142EBFBC7EB8005B55A85B555EF095F50578085BE8FC",
INIT_28 => X"BEAE3D542A004380124921D20975FFAAA1521FF492BF8F40B6AAB84AF555168A",
INIT_29 => X"8F6DE05B40480557A95A3A1C2EBAE28168ABAA2D43D568BC5400168E90E2F412",
INIT_2A => X"47B50A80095178157FEFA0742FA3AA28EA8168A954100071D2E90A855C7A00A3",
INIT_2B => X"0A8F57F6DA971F8F7FFFA42D16D1EAE925EA0BFEBF4AA09217F4905684170851",
INIT_2C => X"000000000000000000000000000002D57AAA8402A8743DBD202DA95568A95E80",
INIT_2D => X"17D34ABA5D7BEAAAAD786BCEAAFFD1564BA2282BFA02A2C28000000000000000",
INIT_2E => X"007F8B2B2D97D483AFA7BD9F5EFA87F57555AAFBD7555FFAE95408A8FDC31AD0",
INIT_2F => X"0A6AEA8FAF0451CA001D4845C2087383F79A5046A37B55F38415555797D63BFF",
INIT_30 => X"A7D7463CC508D07577BAFBD542000D382964A92B401E71D7581C33172EC0A030",
INIT_31 => X"0502828811FCD4EABDB1DFDFC8365A2FD5E04AA5780A8AAAD7AC3CA02003BEBB",
INIT_32 => X"4FF72AAADF245595157050790621F562B1122DA70C3808458881056A5502AA15",
INIT_33 => X"F6A03D4BFB79AFA4C5CB5F5896D55BBAAC55EAFAF86D35E4A92B4460D1506037",
INIT_34 => X"FC0000007FC0000007FC0000007FC0000007FC0000007FC07AAF12E00505D3FD",
INIT_35 => X"7FC0000007FC0000007FC0000007FC0000007FC0000007FC0000007FC0000007",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000400000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"650C00000848A0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000004208B00200E010800006667BE7000102C00080000040012010000080C",
INIT_05 => X"0080000000002020600100208D04414000800000000200004800080000800200",
INIT_06 => X"04022140220932C2038900000100000008082010000000800488000000020400",
INIT_07 => X"088C0060242183060CF118011281B00000220010400020002081A00082100001",
INIT_08 => X"40000400014812466427040098C000622AAAA43E3060C158AC97F0356BDBFBD0",
INIT_09 => X"00026C000559102400200281400469000008B0800000901080004004308B4340",
INIT_0A => X"045413002200000000400408200000201041000208000040020820034200005C",
INIT_0B => X"41E11C008089540000420100101088400000808404004000000020A000100414",
INIT_0C => X"18C191AC191A4191A4191AC191AC191A4191A00C8560C8D08400000609010100",
INIT_0D => X"0E08A20BC417C16004C0B8382210904018000080100100012200000064064019",
INIT_0E => X"0E0615C96000000010200000802100022008100408020401020040100142200E",
INIT_0F => X"C06100000021E300B000000781E00140018000000781E00140018000002430E3",
INIT_10 => X"68C381C00000024E0000000781E00140018000000781E0014001908400005E11",
INIT_11 => X"088400003C30F00C000000155800D00000003E21C0700000000F001180000004",
INIT_12 => X"4000260640900004A400081401A0000004041218503E40300600000048043180",
INIT_13 => X"00009A0001208C30800025200003D807E0000000007252016000904618400013",
INIT_14 => X"480160000F00C0E06100000012D2005100409520381C00000005920004C0C812",
INIT_15 => X"0004025000120850B8180625400400000010711200510004B414780400000055",
INIT_16 => X"1004010040002002080000000804000A0000000011A000100208C008611430A0",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"5800050008000000000000000001004010040100401004010040100401004010",
INIT_1A => X"1451451451564090C69606492492C09A8C205148D757DF8A94102E0001063A29",
INIT_1B => X"BADD6EB75BADD6EB75BADD555555555555555555555555555555555555555145",
INIT_1C => X"FFE0000174BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974",
INIT_1D => X"F5D2AAAB555555400000000000000000000000000000000000000000000303FF",
INIT_1E => X"EFA2D17DEBAF7D1574BAAAFBFDFFFA2FFD74000855555FFFFFFC01FF087BE8BF",
INIT_1F => X"145557BFDEAA5500154AAAAAEBFF455D04175FF5D7FEAAAA002ABDEAA5D2EBFF",
INIT_20 => X"20BAAAD540145F7D5574BAAA8415400005540155F7D16AB45002EA8ABA005540",
INIT_21 => X"975EFF7AEBFF550055555FF55003DE00A2FFFFFEFAAD57DE00082AAAA00082A8",
INIT_22 => X"16AABAAAAEBFE10AAFBD7545F7D5554AA5D2ABDEBA082A821455D2EA8B455D2A",
INIT_23 => X"FFEABEFA2FBEAB455D7BD55FFFF84155FFFFFFFFF55AAAABFFFF5D556AB45A2D",
INIT_24 => X"000000000000175FFF7D140010FF84174BA552EBDEBA0004020AA5D04155FFAA",
INIT_25 => X"4BFBC51FF1471E8BEF55242FF47015A800000000000000000000000000000000",
INIT_26 => X"0B6AEBAEAA5D2EBDFFFBED17FEAAF7D5524AAA2F0BAF7FABDFC7E10005F525D7",
INIT_27 => X"55142A8708202FBD257F1C7550492490E17EAAA2AAB8F4515043DFC75575C700",
INIT_28 => X"03D1420AD000B420820AAE2DB6FB6DF7DFD5038ABA140A2D00554517DEBDB6FB",
INIT_29 => X"25555F8FFDE38087FC51C7F7AABFF55BC5B555C74B8A38E38085BE8B47A3A005",
INIT_2A => X"BA4AF555168B68FEDF6AB52AAABD21EF1C2FEA5FDEBDB505FA4920AFE10082E9",
INIT_2B => X"17AEB8BFF155552B6F5E8BFF1EFBFDBFF5FF1C00BF5D25475C7B7FEAFF45BEAA",
INIT_2C => X"00000000000000000000000000000151EAE3D542A004380124921D20BFFFA0AA",
INIT_2D => X"3D795000087BC01458AFBC11FF55516ABEFDD003EFE5093DC000000000000000",
INIT_2E => X"550434D555C53E0CE2AAA8742BA5D2ABDFFFF7D57DEAAFFD5420B2A2D37DB07A",
INIT_2F => X"F0851575FFAAFBDD5542B2EDD608897FD610D01151C610592A974BAFBAC28B55",
INIT_30 => X"100F3D68FFFAABAC20EF04003FE102400144ABAAFFF7DE772FDD56588042F72E",
INIT_31 => X"4EA0006BFE007E2E8315DD02F6A81A239501755F504BDF557D79431FD006EABA",
INIT_32 => X"03158517BD745AEAEA8FAF0C55EAF57FF957CAAA7FABF7DFD0C6A7DFFFA07FC0",
INIT_33 => X"964A92B403EE18D5408A6F2AFADF6900FFFF68BEFDFFB4B1FE5551141E78A028",
INIT_34 => X"0000000000000000000000000000000000000000000000165BAFBD542000D382",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000400000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0812",
INIT_01 => X"2145A00A1079284D04A044A54E504368404000720885800802000006ECD10200",
INIT_02 => X"5C010800020408040C415854AA055254090541A111000A104A00000009083510",
INIT_03 => X"0C1000100C0000D40526480250149120031500A0218808002440804288890550",
INIT_04 => X"8840C28120051400582012021808040409C0B26850488419444010C10A024A49",
INIT_05 => X"488510910548012025C0C0000300086854B141042252142042A048D090006372",
INIT_06 => X"948037480159A403109848000428AA8282102040449090D520085224410AA420",
INIT_07 => X"01020402242000408468112010810C055200022025A83AA3008882004A001542",
INIT_08 => X"11491C154429220A2824640010A010020282843E0008124C0000211000008840",
INIT_09 => X"E280442C1411D020828A2B116824632885419240016001900AE01A2020066395",
INIT_0A => X"30105108880684145002021012D40D718241108815380200900160AE42CE2818",
INIT_0B => X"53419F10308D100054AA080092112C100B400880454058E80B94080C49318000",
INIT_0C => X"D0090D0090D2890D0890D2890D0890D2090D0048610486808403A384880B8981",
INIT_0D => X"8202043800000620500403080A919000B8AD0304144008111A00582043243050",
INIT_0E => X"9835300002AA40AA902408200010002021060C810241832241280C81A0984020",
INIT_0F => X"100000000080A0000140000002000140200A8000000200014020100290E469C6",
INIT_10 => X"00100000000003400A8000000200014020094000000200014020087000000000",
INIT_11 => X"014200000004000000000081400004C00000000020000000008C000010A00000",
INIT_12 => X"0510000000000006800001880004008400800000000020000000000048100000",
INIT_13 => X"0000D0260000000000003409280000000000000040025000030000000000001A",
INIT_14 => X"400002A0000000000000000042900000A100000000000000008012A200000000",
INIT_15 => X"000000004420300000000000000000000010C010000098000000000000000105",
INIT_16 => X"00802208036408C0820010004D36A222120090554000E40080000000088000A0",
INIT_17 => X"8802008020080200822088220882208802008020080200822088220882208802",
INIT_18 => X"8320883200812008120081208832088320883200812008120082208822088220",
INIT_19 => X"E88051029FC0FC0FC1F81F81F820883208832088320081200812008120883208",
INIT_1A => X"08208208208C13A4301040B2CB2CBAC838B6C0080271AE180616A851158E2863",
INIT_1B => X"944A25128944A25128944A082082082082082082082082082082082082082082",
INIT_1C => X"FFE381F928944A25128944A25128944A25128944A25128944A25128944A25128",
INIT_1D => X"A550002000AA800000000000000000000000000000000000000000000003C200",
INIT_1E => X"BAFFAE801FF087BE8BFF5D7BEAA1055042AA105555421EFFFD568AAA002EBFEB",
INIT_1F => X"FFFA2D57DE10557BE8ABAF7AAA8BEFAAAE975FFA2D5555450851574000851554",
INIT_20 => X"5555F7D568ABAF7D5574BA552EA8AAA5D2EBFFFFA2D1554BAF7D17FEBAAAFFFD",
INIT_21 => X"EAAAA552AAAAAAAAAABFF455D04175FFFFD5574AAAAAA974BA082EA8BEFAAD55",
INIT_22 => X"FEAA000055401555D7BFFE10085557410F7AA97410087BD55FF087FEAA10A2FF",
INIT_23 => X"0017400550402155A2803FE005D7FE8B45F7FBFDE00085540155F7D56AA00007",
INIT_24 => X"00000000000017400082AAAA00082A820BAAAD540145F7D557410AA8428A1055",
INIT_25 => X"4BD16FAAA002ABFEAA550E82000E28A800000000000000000000000000000000",
INIT_26 => X"FEAFBD2410005F57482E3AA801FF1471E8BEF5574AFA00010ABFA38555F401D7",
INIT_27 => X"AAF7D5524AAA2F1FAF7FABFBFF400417FEF082F7AAA8BEFE2AA955EFA2DB5757",
INIT_28 => X"492082EADBFFBEDB55555E3DF6DA82F7DF520385D2FE80AA5D2EBDFD7BED1574",
INIT_29 => X"21C7005B6FB47F7A438E925D24ADAAAB6AAB8F455784155C75575C7000B6AE95",
INIT_2A => X"4717DEBDB6FA3D0075EDA800051C05571474024A81C5557578EBA087400007FC",
INIT_2B => X"FFDE381D716FA15550015428E10A001FFB40038F68F7F578F7FFEF568E280855",
INIT_2C => X"000000000000000000000000000001043D1420AD000B420820AAE2DB4716DF7D",
INIT_2D => X"828FDEBA5D7BC015582D57DEAA002ABDEAA552A80010AAA88000000000000000",
INIT_2E => X"AAAE955EFAAFBC15F5A3D7D6800087BD5410AAAA801FF55556ABEF5D517EEE00",
INIT_2F => X"A5D2ABDF55F7D575EAAFFD50A2B2A3D169B07A3D7BFE10597BFDE00AEAC28BFF",
INIT_30 => X"555A53C00B2A2AA02000082ABDFEFFFFBC1154AAFFFFE107FF9D72A20842080B",
INIT_31 => X"4EAA28015400547FC315D00797CF4780286A2105D2A3FEBAFFAC28B555504145",
INIT_32 => X"99ADABD5A8AAA0051575FFA2FFFDA02003FFDEAA8557D65550915544AA5D5157",
INIT_33 => X"144ABAAFFD75E7F2BDDD2B8016F9E2555500174AA282E20BFFFF842AAAAADD56",
INIT_34 => X"0000000000000000000000000000000000000000000000030EF04003FE102400",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000800000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380206",
INIT_01 => X"200C9A40408001683C0462C99E004B61404040028804A0080A000416A0990A0C",
INIT_02 => X"4809A900031800444461089866E331352180D468B8040E600C0081110B802CD0",
INIT_03 => X"6D0B61108C00014231A3080408C68420330066010A80881068A808401CC46330",
INIT_04 => X"482218066A09C03B348C1C1928DD5A4402211A68470944842640902107002D24",
INIT_05 => X"0583180353202020000144E50B44644B30A86D05014A0D224063095092100E34",
INIT_06 => X"54023740216934020303680A040066D98A182210085A50C02048288234629414",
INIT_07 => X"018C00220430814204E01C581291820CCA000E3226413990008C80205A00CCCC",
INIT_08 => X"4108747320081246252D5010184000220002A43E10294258E805E1156002D940",
INIT_09 => X"D0AA546AC41B112029A61D84424429AA1320B1010140C1350B48292020024180",
INIT_0A => X"000102022850A1CC0047071913208CE802430488082042008040F399606F4058",
INIT_0B => X"5141BE42B88840005268081412152900484201A814144D60888CAA2C48151020",
INIT_0C => X"1B49019490194901B4901B4901949019C901B64805E480CA94480506980125C4",
INIT_0D => X"5A01E2B1080602E00C54216800859000199C98800C8140A11A44423040240450",
INIT_0E => X"28A65300E6664599902600009821204A040C1C040C0205038300480801480208",
INIT_0F => X"000000000090000003202900000010002008A02900000010002008039666928B",
INIT_10 => X"00000000000801000A202900000010002009E0290000001000200A3800008000",
INIT_11 => X"036000008000000000000088000002D003008000000000000280100016200812",
INIT_12 => X"05B008088000008201021C880000488002810005000000000000040000100000",
INIT_13 => X"0010402B80412000000410199800040000000000408020000680209000000208",
INIT_14 => X"800012980040300000000000C020000C8300208800000000008200AE01011000",
INIT_15 => X"40A0000841003100010401000000000002008020000C38000200000000000120",
INIT_16 => X"10070300704028820801400068360424820185CCE0128010020000008088021C",
INIT_17 => X"0070100701007010050180501805018050180501805018070100701007010070",
INIT_18 => X"070140601007014060100701C040180501C040180501C0401807010070100701",
INIT_19 => X"4A81454A26AA555AAB554AAB5541C040180501C040180501C040180501406010",
INIT_1A => X"08208208209441D0B0000092492480AA2860607818F18E0C851428200B262C31",
INIT_1B => X"D4EA753A9D4EA753A9D4EA492492492492492492492492492492492492492082",
INIT_1C => X"FFD55E21A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8",
INIT_1D => X"FAA8000155080000000000000000000000000000000000000000000000000200",
INIT_1E => X"EFFFD568AAA002EBFEBA555142000AA802AA10F7D57FEAA557BE8B45A2D5555E",
INIT_1F => X"A10550402000AAD56AAAA557BC0155A280021EFA2FFE8B4555042AA105555421",
INIT_20 => X"0010AA842AAAAFFD542000FFD5574000851554AAFFAE801FF087BC01FF5D7FEA",
INIT_21 => X"7DE105551420BAF7AAA8BEFAAAE975FF005540145A2D157410AAD17DFFF5D040",
INIT_22 => X"03DEBAAAFFFDFEFAAD57DEAAF7AE975FF080428B455D7FFDEAA5D55574BA0051",
INIT_23 => X"AE800AA087BD5555552A821EF007FFFEAAAAD5554AA552EBFFFFA2D5554BAF78",
INIT_24 => X"000000000000020BA082EA8BEFAAD555555F7D568ABAF7D5574BA552E800BAAA",
INIT_25 => X"E975EAB6DBEDF575FFAA8E02155080E800000000000000000000000000000000",
INIT_26 => X"5EBAEADA38555F451D7EBD16FAAA002ABFEAA555E02000E28AA8A38EBD578E82",
INIT_27 => X"FF1471E8BEF5575EFA00012A87A38AAD56DA824975C217DAA84021FFAAF5EAB5",
INIT_28 => X"400BED57FFD7410E05038BE8E2DABAFFDB47412ABFE90410005F57482E3AA801",
INIT_29 => X"FEBA5D71D742A407FFFE00555F47082E3AAA8BEFA02A955EFA2DB5757FEAFBD2",
INIT_2A => X"BFFD7BED157482F7803AEAAA2F1FAF7FABFBEAE2AEBA4974871C043AB6D4975F",
INIT_2B => X"F7AE38497FC00BAB6A4850821C75D25C74920821D708757AE2AA3FFC04AA552E",
INIT_2C => X"0000000000000000000000000000007092082EADBFFBEDB55555E3DF6DA82F7D",
INIT_2D => X"AA8A8ABAAAD568A1020516ABFFFFFFD75FFAAAE8014500288000000000000000",
INIT_2E => X"AA80001FFAAD57EB55A2A8ABEBA5D7BD5545A2D57DEAA002EBDEAA557BC0010A",
INIT_2F => X"0087BD5410AAAA801FF5555629EF5C517EEE00828D74AAFBD57DE000057C21FF",
INIT_30 => X"EFA8FBC15E5A3D5D7400FFD57DF55082E974AAFFAABDEBA77FDD66A0ABBDC200",
INIT_31 => X"50555002ABFF54517EEB25D57C14100957FF6105D7BD5400AAAC28BFFAAAE955",
INIT_32 => X"FA42A3D7020BA5D2ABDF55F7D1554A8FFC42AA10A7D169F57ABD7FEEBAAA8415",
INIT_33 => X"C1154AAFFFFE10FFF9DF202096F014AAFF84154105555C215500000014558557",
INIT_34 => X"000000000000000000000000000000000000000000000015400082ABDFEFFFFB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000400000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204002",
INIT_01 => X"01039802000820491C00650E1E004340403008418984014902030906A8D10200",
INIT_02 => X"480108A000000000444048E41E80F00A41043118680002000800000009882390",
INIT_03 => X"06504110080000D0040608024010102026001260300000003080880208C000F0",
INIT_04 => X"9100E98268154C1AE0B01C160033B944028290285AE0DC38E02090E81C22E801",
INIT_05 => X"5C0F20B36F000109200044C401041C4CF21C48B433483C8242EAE1B0000074C4",
INIT_06 => X"100007000059800310086A1A0022E18780000140C9D9D0930000F228075A6071",
INIT_07 => X"00000000242000008461000810818403C100060064012E00048C82201800BC28",
INIT_08 => X"0048CC8F01090602202C0400008000002202243E400010480000211540008810",
INIT_09 => X"40E0DC1EB5191120C7BE7D152201612E80E891E0614041340838450020422111",
INIT_0A => X"30545DAD8C2E0982400603003200872003FB1408082840002044007846164E0A",
INIT_0B => X"43411D10118D1A04522E000498140C104B260DA0404003C08B6000AC01128000",
INIT_0C => X"C5010C3010C1010C3010C1010C1010C3010C140869808618850BE6305989AB80",
INIT_0D => X"100140302800108018840440028480001B8780800000003102045C3443043410",
INIT_0E => X"3080620481E0E18790012A001001026808000002020101028100200180080201",
INIT_0F => X"000000000010000005C0200000001000000C4020000000100000000380E4C308",
INIT_10 => X"00000000000800000D00200000001000000EC020000000100000086A20008000",
INIT_11 => X"012820008000000000000008000001B00100000000000000020000002AA00010",
INIT_12 => X"06D0000080000080000241D80000800442800001000000000000040000000000",
INIT_13 => X"0010003A00002000000400021800040000000000008010000B00001000000200",
INIT_14 => X"400005900000100000000000801000089000008000000000000200F800001000",
INIT_15 => X"00000000A500100000000100000000000200001000002E000200000000000020",
INIT_16 => X"000000C032700000022400444934240A8021B63C005108010004100098098010",
INIT_17 => X"C010080200401008000040300800004010000200C01000020040100802004030",
INIT_18 => X"02000000000100C0300400008000000300C0100C00000020080000C030000000",
INIT_19 => X"20240142325930C9A6CB261934C000200801004030040200800000030040100C",
INIT_1A => X"14514514514E98264686668A28A260521CC45140C700FC0A0002870980831A28",
INIT_1B => X"1A8D46A351A8D46A351A8D555555555555555555555555555555555555555145",
INIT_1C => X"FFD5E7D8341A0D068341A0D068341A0D068341A0D068341A0D068341A0D06834",
INIT_1D => X"A5D55420AA002A80000000000000000000000000000000000000000000000200",
INIT_1E => X"AA557BE8B45A2D5555EFAAD140155080000155FF843FFEFAA84001FF5D043FEA",
INIT_1F => X"000AA80001555D04174AA002A80010FFAE975FFAA80001EFA2AAAAA10F7D57FE",
INIT_20 => X"00BA5D51555EF002AA8BFFAAAAAAA105555421EFFFD568AAA002EBFEBA555542",
INIT_21 => X"82000AAD568AAA557BC0155A280021EFA2FFE8B45F78400145FF842AAAAA2AA8",
INIT_22 => X"BC01FF5D7FEAA105D0428B4500003DFEF080428B455D002AABA5D2AAAAAA5D2E",
INIT_23 => X"80154BAA2FBE8AAAF7AA821EFAAAAA8BEF552E820000851554AAFFAA801FF087",
INIT_24 => X"00000000000015410AAD17DFFF5D0400010AA842AAAAFFD542000FFD57DF55A2",
INIT_25 => X"A284051D755003DE92415F42092142E000000000000000000000000000000000",
INIT_26 => X"71C0A28A38EBD57DE824975EAB6DBEDF575FFAADE02155080E85145E3803FFEF",
INIT_27 => X"AA002ABFEAA555F42000E2AA851455D0A124BA002080010FFA4955C7BE8E021C",
INIT_28 => X"145F7802AABAA2A480092415B505D71424AABD7F68E2FA38555F451D7EBD16FA",
INIT_29 => X"AA824924AAA92550A07038BED56DA824975C217DAA84021FFAAF5EAB55EBAE82",
INIT_2A => X"55482E3AA801FF1471C01EF5575EFA00012ABFB6D080A3AFEF080A2FB45490E2",
INIT_2B => X"B6FA12ABAEBDF7DAA80104BAAAFFEAA00F7AE821D7B6A02FBC71D0E10010005F",
INIT_2C => X"0000000000000000000000000000010400BED57FFD7410E05038BE8E2DABAFFD",
INIT_2D => X"02897555A2803FFFFAA841754555043FE10087BC2000552C8000000000000000",
INIT_2E => X"FF8017545F7AE821455D2CAAABAAAD57DE1000516ABFFFFFBD75FFAAFFC01450",
INIT_2F => X"A5D7BD5545A2D57DEAA002EBDEAA557BC0010AAA895555042E820BA080400010",
INIT_30 => X"FFAAD57EB55A2A880155F7802AAAAAA8002010007FC0155D5022A955FFACBFEB",
INIT_31 => X"BEF002EBDF45542AAAA0008043CAB0552C97CAAFFD57DE000057C21FFAA80001",
INIT_32 => X"CFE55D2CC2000087BD5410AAAA801FF5555421EF58517EAB00028A9BEF002EAA",
INIT_33 => X"974AAFFAABDEBAF7FDDE6A0AA90FDFEFA280020BAA2FFEAA10FFAE82145F7803",
INIT_34 => X"000000000000000000000000000000000000000000000002000FFD57DF55082E",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000800000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A337A20E07C0C1E006",
INIT_01 => X"295FBC468000A04D5C6A60000C34C24841280A00084000C8C212892EEAD53235",
INIT_02 => X"C809AD5CB118E640A4D158F8011FF0002080000082C8C66609DB7DDDCB1F2036",
INIT_03 => X"250906263A4C904214A35C80085285720B20648A88800000B8E0F852A884500E",
INIT_04 => X"4005122126899100064D20001044429C78A43A2C4436CC87198A3916E0551A24",
INIT_05 => X"A370C14CA0E900004048402389CFE2F20F7D7A354CB5C208E51437F044948912",
INIT_06 => X"9B9407B9424F33468B096FCF452AE0505A185905CC2414D44437118630839B88",
INIT_07 => X"588C732074A68D5AB4EB180717FF513FC52691924098712CE481FDC201D43C1A",
INIT_08 => X"0016053F180A1286A4ED1BC18840C320000055FE91AA545CBA4DE1D17992D9BE",
INIT_09 => X"2D1A4D8105B734723041008100486100601EDE1DE46431138DFD404CB4022595",
INIT_0A => X"A131112C0D15C901B2122309204C28B67061E81A8920C8D3CF8014007902DA6B",
INIT_0B => X"AD5C3402488888E5126BA350B27C092E63D18C9C500577EEA33EF24C09B42464",
INIT_0C => X"096B80D6B80B6B80F6B8096B80F6B80B6B80D15C04B5C07AD50C94020D233107",
INIT_0D => X"8948020D829FA454104132252011E542387F810480C840C383751EF5606E0178",
INIT_0E => X"000200CA7FE0627FD25845E42151648F854480A042512028100A8C38280AA04C",
INIT_0F => X"D06101C55DE5E3E3C017E37FC3E0017C3F8817E37FC3E0017C3F900040241001",
INIT_10 => X"6CD381C0118797FE0817EA7FC3E0017C3F8817EA7FC3E0017C3F9900DFFFDE15",
INIT_11 => X"F800DFFFBE34F00C0270F3F55F1F8007FDBEBE25E0700463E1FF2C7E014FF7BE",
INIT_12 => X"C5DEF64EC090626FE40140459759173BBD6EF37D523E6030061341F07FD571F8",
INIT_13 => X"0C4DFE2A6FE2AC3082637F281BFFFC07E00007E07F7253D38337D1D6184131BF",
INIT_14 => X"4F4F8397FFA0F0E06101C53E76D3D3E884FDDDA8381C0098E5FD92BBDFC8D812",
INIT_15 => X"19074FA36FDF58DBF81C072540049707E0FEF313D3E03BFFF61478040570EFD5",
INIT_16 => X"8CA02ACA00C50850182309444D248204201040FC190054A2110B8ACC483204A1",
INIT_17 => X"0A128CA0284A2280A1288A128CA2284A0288A1288A3284A228CA0288A1280A32",
INIT_18 => X"A228CA0284A3280A3288A1288A3280A2284A028CA2284A2284A028CA0280A328",
INIT_19 => X"F6A1850E1892596D34924B2DA6A84A2284A1288A1280A3280A1288A0284A2284",
INIT_1A => X"7DF7DF7DF7CBFBFE7EFEEE79E79EFAF3F51EB769CFEF73B6FFE74FC2400DB6DB",
INIT_1B => X"EEF77BBDDEEF77BBDDEEF77DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF",
INIT_1C => X"FFC27F6BDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDD",
INIT_1D => X"55D2E955FFF7FFC0000000000000000000000000000000000000000000000200",
INIT_1E => X"EFAA84001FF5D043FEAA5D04020AA002AAAABA555140155087FFFFEF00042AB5",
INIT_1F => X"1550800001FF5D00001555D2E975FF5D5568B555D7BD5545FFD540155FF843FF",
INIT_20 => X"FF45A2FFC0000AAAE974AAFFFFEAA10F7D57FEAA557BE8B45A2D5555EFAAD540",
INIT_21 => X"401555D04174AA002A80010FFAE975FFAA80001EF002AAAABAF7D168A10A2D17",
INIT_22 => X"EBFEBA555542000A28028BFFF7803DF55FFAEBFE005D2EAAB45557BD55555555",
INIT_23 => X"517DF55082E974BA087FE8B55552E955EF5D7FEAA105555421EFFFD568AAA002",
INIT_24 => X"00000000000000145FF842AAAAA2AA800BA5D51555EF002AA8BFFAAAA820AA5D",
INIT_25 => X"007FFFFFF1C042FB7D492A955C7F7FBC00000000000000000000000000000000",
INIT_26 => X"5E3DB45145E3803AFEFA284051D755003DE92410F42092142E28ABA5D5B4516D",
INIT_27 => X"6DBEDF575FFAADF42155082E851C75D0E02145492E955C75D5F6DB55497BD554",
INIT_28 => X"ABAF7D16DA28A2DB7AF7DB6FBC7028A2AA95492FFFFE8A38EBD57DE824975EAB",
INIT_29 => X"FB45557BD5555415F45145490A124BA002080010FFA4955C7BE8E021C71C0A2D",
INIT_2A => X"451D7EBD16FAAA002ABFEAA555F42000E2AAA8BEFE3843AF55E3AABFE105520A",
INIT_2B => X"4821D7F68E07082495B7FF7D082E954AA087FEDB7D5D2A155D7157BEFA38555F",
INIT_2C => X"0000000000000000000000000000002145F7802AABAA2A480092415B505D7142",
INIT_2D => X"52CAAAAA5D7FD75EF087BFDFEF5D003DFEF002E95555F7FDC000000000000000",
INIT_2E => X"5D7BFDF45007FD7555A2F9D5555A2802ABFFAA841754555043FE10082A820005",
INIT_2F => X"AAAD57DE1000516ABFFFFFBD75FFAAFFC0145002895545552E80145002E95545",
INIT_30 => X"45F7AE821455D2CBFEAAFFD17FEAAAAFFEABFFF7FFD54BAA2AA95410F7FDEAAB",
INIT_31 => X"B45AAAABFE0009043FF555D7BD55550879D5555002E820BA080400010FF80175",
INIT_32 => X"75455D7DFFEBA5D7BD5545A2D57DEAA002EBDEAA557BC0000AAA8A8BEFA28028",
INIT_33 => X"02010007FC0155550222955FFAC97400087FFFFFF002E954AA087BFFFFF5D2E9",
INIT_34 => X"000000000000000000000000000000000000000000000000155F7802AAAAAA80",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000003000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B0061A258A2840112C03002C180004003220200403302301C0381A0086",
INIT_01 => X"860041C83839484C00A100000052024841000000090800090210010000510204",
INIT_02 => X"080108200C1000004464080400C0080100000000010432400800800009882050",
INIT_03 => X"040001008C2340D0800208624200002183800584488000103080010C08C10000",
INIT_04 => X"00101610A029B08400044800000000040008102A040810040400900500001800",
INIT_05 => X"02800000400C830934E4A0002900404400820000000A00824004084011200A00",
INIT_06 => X"14C8874C884D0C024608680210C11F8010122100880802800308010000829400",
INIT_07 => X"060800002430200004611000508184803A0900224000200008818028C04883E1",
INIT_08 => X"4041FE80E009024260240010608000000000043E040000488000201400008810",
INIT_09 => X"0002447E041B112020208010404029006FE0B081003204502000002068621191",
INIT_0A => X"35E5148B0D916BBE39049191200000200441048108000220002FC5FA60000148",
INIT_0B => X"5358BF12E88D1000022808801A112D1443142A815440600083FE9AA300100281",
INIT_0C => X"C1416C1416C5416C5416C3416C3416C7416C500B60A0B60AD40E34104C093904",
INIT_0D => X"8C03403C440C054048850A300A8480009A0020865AE4ECB11B441A105B05B016",
INIT_0E => X"00000031001E4800022100321489214001A742D3A368D1B4686D100234B44242",
INIT_0F => X"00000000000AB800302008000000014000602008000000014000674000260000",
INIT_10 => X"0000000000000241E020010000000140006020010000000140006A8400000000",
INIT_11 => X"028400000000000000000003C00052000200000000000000000CD00184000800",
INIT_12 => X"30000800000000049A48184000A0400000010000000000000000000048028C00",
INIT_13 => X"0000918480010000000024C9E000000000000000000FF0006440200000000012",
INIT_14 => X"C000602800400000000000000BB000112B0020000000000000007E0000010000",
INIT_15 => X"02A0005000202500010000000000000000104CF000198000000000000000000F",
INIT_16 => X"4AD2B46D180684E8402440044C24A30819020603E0A20640C8400010218432A0",
INIT_17 => X"2D1B4ED3B4AD0B42D1B4ED2B42D0B46D1B4ED2B42D1B46D3B4AD2B42D1B46D2B",
INIT_18 => X"D1B42D0B46D2B4AD1B46D0B4AD3B4ED0B46D1B4AD2B4ED1B42D0B4ED3B4ED0B4",
INIT_19 => X"F8840000331C618E38E38C31C7346D3B4AD3B46D0B42D3B4ED2B42D1B42D2B4E",
INIT_1A => X"1C71C71C71CEDBB676F66EFBEFBEFAF99CFEF179CFF1FE1E9F52AFF9BFAFBE7B",
INIT_1B => X"FE7F3F9FCFE7F3F9FCFE7F1C71C71C71C71C71C71C71C71C71C71C71C71C71C7",
INIT_1C => X"FFE43591FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"05D2EBDF55557FC0000000000000000000000000000000000000000000030200",
INIT_1E => X"55087FFFFEF00042AB555D2E955FFF7FFC21EFF7D17DEAA5D2AAAAAA5D557DE1",
INIT_1F => X"0AA002A82145555542010FF803DEAA5D5568BEF5D042AA10A2AAAAABA5551401",
INIT_20 => X"20BA00557DF455D7BFFEAA555540155FF843FFEFAA84001FF5D043FEAA5D0002",
INIT_21 => X"001FF5D00001555D2E975FF5D5568B555D7BD5545FFD568AAA5D00154AAAAD14",
INIT_22 => X"5555EFAAD540155080000000F7843FF55007FFDEAAA284020BAAAD168BFF0800",
INIT_23 => X"51401EFF7842AA00FF8417545AAAEBFE10FFFFEAA10F7D57FEAA557BE8B45A2D",
INIT_24 => X"0000000000002AABAF7D168A10A2D17FF45A2FFC0000AAAE974AAFFFFC21EF55",
INIT_25 => X"5520ADA92495B7AE10412EBFF45497FC00000000000000000000000000000000",
INIT_26 => X"0AAAAA8ABA5D5B4516D007FFFFFF1C042FB7D492A955C7F7FBC71EFFFD57FE82",
INIT_27 => X"D755003DE92410E02092140E0716D415F47000F78A3DE92415F6ABD7490A28A1",
INIT_28 => X"A92550A104AABED1470AA005F78F7D497FFFE925D5B45145E3803AFEFA284051",
INIT_29 => X"20BAA2DB68BC7140E051C75D0E02145492E955C75D5F6DB55497BD5545E3DB6A",
INIT_2A => X"7DE824975EAB6DBEDF575FFAADF42155082E87038FF8038F6D1C7BF8EAAAA800",
INIT_2B => X"A95492FFFFC71EF415F471C7FF8428A00E38412545AAAE3FE10A3FBE8A38EBD5",
INIT_2C => X"000000000000000000000000000002DABAF7D16DA28A2DB7AF7DB6FBC7028A2A",
INIT_2D => X"7FDD55EFF7D57DE005D003DE00007FEAA10002ABFF450079C000000000000000",
INIT_2E => X"087BE8B45082EAAA10A2A8AAAAA5D7FD75EF087BFDFEF5D003DFEF002E95555F",
INIT_2F => X"5A2802ABFFAA841754555043FE10082A82000552C955FF007BD5410FFAABFE00",
INIT_30 => X"45007FD7555A2F9EAA005D2A820AAF7D5574AA087BEABEF007FFDE00557DD555",
INIT_31 => X"BFF557BE8ABAA284020BAA2FBEAB55552C95545552E80145002E955455D7BFDF",
INIT_32 => X"FE10A2F9EAABAAAD57DE1000516ABFFFFFBD75FFAAFFC01450028974BAFF842A",
INIT_33 => X"EABFFF7FFD54BAA2AA95410F7FDD55EF007BD5555F7802AA10AA8000145AAAEB",
INIT_34 => X"00000000000000000000000000000000000000000000003FEAAFFD17FEAAAAFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000002400000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0048201002842002C02450018800002300500030B313300C418992002",
INIT_01 => X"A34009C23838684D1C20E0000E11426840000000080000080200080000110200",
INIT_02 => X"4801082048100000446558040080000041000000000622400800000009000010",
INIT_03 => X"040001818CA144D0842248424210812103000480088000003080014688800000",
INIT_04 => X"000012002041900000048000000000040088322944200C850001940400301800",
INIT_05 => X"0200000040084000284000204104004402000025000800065004207030320800",
INIT_06 => X"108017080149000246086A2A1468004012120004440812D40120008200829001",
INIT_07 => X"2408000024302040846810005281848003494020400031240C8C8218E06A0009",
INIT_08 => X"4040050001090242602C0418408000000000243E0408104C8000201540008810",
INIT_09 => X"00024401041B132820000001424069004000B204636009104A0101226A422104",
INIT_0A => X"80049800A0281400300B0210200008B206639389480046240068180262000048",
INIT_0B => X"41401C1081811C44D22A18841616004118004482040448011800004D49340082",
INIT_0C => X"00192001920019200192041920419204192060C9010C90100008040008012101",
INIT_0D => X"48A000880144434A001001228000803198003604004048294008C40C483480D2",
INIT_0E => X"0000002160006000100000200811020805000480004000220108000060000800",
INIT_0F => X"09864038A2881210382000000001E003E0582000000001E003E0422834240000",
INIT_10 => X"0000160700706901982000000001E003E0582000000001E003E04E8400000000",
INIT_11 => X"0684000000000330C00F0C8210807200000000000581C01C1C809201C4000000",
INIT_12 => X"29D000000C2419121028C00020A2400000000000080082C180603A0E003A0904",
INIT_13 => X"8322414E800000432118908DF8000000061E001FC00C10207740000021908C48",
INIT_14 => X"40806BB800000009864038C14810201BAB000000026130071A80613A00000184",
INIT_15 => X"840080546520350000600812058100F81C018890201BBA0000008239020F1108",
INIT_16 => X"04812208033400C0022140404D268624B210040004A08400000044222900320C",
INIT_17 => X"0832048120481204822008020080204832048120480200802008020081204812",
INIT_18 => X"802008020C812048020080200812048120080200802048120483200802008020",
INIT_19 => X"0221054A2C208200010410400020880200812048120C80200802008120C81200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFD3B3D800000000000000000000000000000000000000000000000000000000",
INIT_1D => X"5AA8017410555540000000000000000000000000000000000000000000000200",
INIT_1E => X"AA5D2AAAAAA5D557DE105D2EBDF55557FFDE00557BEAABAA2AEAABEFF7801555",
INIT_1F => X"5FFF7FFD5555557BEABFFF7FBEAAAAAAD157555AA803FEBA5555421EFF7D17DE",
INIT_20 => X"DFEFAA80000BAAAAA820BAA2802AABA555140155087FFFFEF00042AB555D2E95",
INIT_21 => X"02145555542010FF803DEAA5D5568BEF5D042AA10A2AA955EFF7FFD5400F7FFF",
INIT_22 => X"43FEAA5D00020AA002ABDEBA5D7FE8A000004154BAF780001EFAAAAA8B450000",
INIT_23 => X"2AAABFF5551421FFAAD157545AAD5555EF557FC0155FF843FFEFAA84001FF5D0",
INIT_24 => X"00000000000028AAA5D00154AAAAD1420BA00557DF455D7BFFEAA5555575455D",
INIT_25 => X"AAA0A8BC7EB8417555AA84104385D55400000000000000000000000000000000",
INIT_26 => X"A4155471EFFFD57FE825520ADA92495B7AE10412EBFF45497FFFE385D71E8AAA",
INIT_27 => X"FF1C042FB7D492A955C7F7FBD056D5D75EABC7FFF5EAAAABEDF5257DAA8438EB",
INIT_28 => X"5EFEBFFD2400EBFBFAFEFAA80070BAA2A0870BAAA8028ABA5D5B4516D007FFFF",
INIT_29 => X"01D7AAA0AFB6D1C040716D415F47000F78A3DE92415F6ABD7490A28A10AAAA92",
INIT_2A => X"3AFEFA284051D755003DE92410E02092140E3DE924171E8A281C0E10482F7840",
INIT_2B => X"FFFE925D5B525454124AFBC74955421EFA2DF5557DAAD5D05EF0175C5145E380",
INIT_2C => X"000000000000000000000000000002AA92550A104AABED1470AA005F78F7D497",
INIT_2D => X"079FFEAA5D5568ABAA2842AB55A28015545A284000BA5D534000000000000000",
INIT_2E => X"F7FBC01EFA2842AABA0857555EFF7D57DE005D003DE00007FEAA10002ABFF450",
INIT_2F => X"A5D7FD75EF087BFDFEF5D003DFEF002E95555F7FDC01EF55556AB55F7D56AABA",
INIT_30 => X"45082EAAA10A2A8801FFA2FFC2000A2FFEABFFAA84174BAAA80174AAAA862AAA",
INIT_31 => X"AAA552A80010F78000145AA843DFEF5D02155FF007BD5410FFAABFE00087BE8B",
INIT_32 => X"21FF085755555A2802ABFFAA841754555043FE10082A82000552CBFE10085168",
INIT_33 => X"574AA087BEABEF007FFDE00557DC014500003FF450051401FFA2FBD55EFAAD54",
INIT_34 => X"00000000000000000000000000000000000000000000002AA005D2A820AAF7D5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"A14008420008204D042100000212026840000000180800080200090048510204",
INIT_02 => X"080108000090000004655C040080000051000000000402400800000009000010",
INIT_03 => X"00000100803008D0842240024210810003800584488000103080894288800000",
INIT_04 => X"00009610A028B084000440C0040000040088323244280C950400808500321800",
INIT_05 => X"42800080400C8A09306420202804400402800035200A00020204287001114A00",
INIT_06 => X"14C8864C8849880002486800142BFF001292214444081254002801A200821400",
INIT_07 => X"004800002430204084281000D281040001182020400031241C0D80000041BFE9",
INIT_08 => X"444005000108020220240010048000000000043E0408104C8000000100008810",
INIT_09 => X"0812040105191100200081130210ED104008A285617205D02A01010141225091",
INIT_0A => X"8004C8252291490039039390200008B20E230008280040088040100240008061",
INIT_0B => X"40013C128BC95C44522A00241204094008442681100448000800826F49240001",
INIT_0C => X"0408000080000800008000080000800008000440020400229548040008012125",
INIT_0D => X"401140BC4028430108150900408590109A00209642E46CA00240460400200440",
INIT_0E => X"080410010000200002210A320C89000005A142D0A16850B6294D100234201242",
INIT_0F => X"2F9EC00000800008100020003C1FE00020080020003C1FE00020044014260082",
INIT_10 => X"132C7E3F00000100080020003C1FE00020080020003C1FE000200880000081EA",
INIT_11 => X"0080000081CB0FF3C000008000201000010001DA1F8FC0000080110080000010",
INIT_12 => X"040000B0BE6C00020040580040200000001004832CC19FCF81E0000000100002",
INIT_13 => X"80004020000C31CF60001000000007F01FFE00004000300420000618E7B00008",
INIT_14 => X"C0102000000F151F9EC0000040300401000200D547E3F00000800080001617AD",
INIT_15 => X"02A020100000822406E1B95A3F83000000008030040100000BAB87FB00000100",
INIT_16 => X"46D1B66D1A368C68D26000544D26A504AB120400222206404840001101843000",
INIT_17 => X"2D1B46D1B46D1B46D1B46D1B46D1B42D0B42D0B42D0B42D0B42D0B42D1B46D1B",
INIT_18 => X"D1B46D1B42D0B42D0B42D0B42D1B46D1B46D1B46D1B42D0B42D0B42D0B42D0B4",
INIT_19 => X"20840442200000000000000000346D1B46D0B42D0B42D0B42D0B42D1B46D1B46",
INIT_1A => X"3CF3CF3CF3DBF91E66C6FAD96D965201F4C251414A87D78AF421448BE28F3AEB",
INIT_1B => X"3E1F0F87C3E1F0F87C3E1F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"FFD160B27C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C",
INIT_1D => X"AFFFFC2000557FC0000000000000000000000000000000000000000000000200",
INIT_1E => X"BAA2AEAABEFF78015555AA80174105555420000000021EFAA843DE00F7803FEB",
INIT_1F => X"F55557FD54AAA2AA955FF00043DE005504175FF08514014555557DE00557BEAA",
INIT_20 => X"DF45FFD17DFFFFFD56AA00557FC21EFF7D17DEAA5D2AAAAAA5D557DE105D2EBD",
INIT_21 => X"55555557BEABFFF7FBEAAAAAAD157555AA803FEBA55556ABFFA280154BAFF803",
INIT_22 => X"42AB555D2E955FFF7FFD5410002AAAAAAA2D57DF450004154BA087BEAAAAF7D5",
INIT_23 => X"843DE1008556AA00A28028B55FFD1555EFA2802AABA555140155087FFFFEF000",
INIT_24 => X"000000000000155EFF7FFD5400F7FFFDFEFAA80000BAAAAA820BAA280000AAA2",
INIT_25 => X"A2803AE38FF843DEBAEBFFC20285D75C00000000000000000000000000000000",
INIT_26 => X"55D5F7FE385D71E8AAAAAA0A8BC7EB8417555AA84104385D5542038000A001C7",
INIT_27 => X"92495B7AE10412EBFF45497FD24BAA2AA955C708003FE285D00155FF00554515",
INIT_28 => X"BEFA28E124AAF7843AF7DEBDB78FFFE3DF6DA284175C71EFFFD57FE825520ADA",
INIT_29 => X"04920875EAA82F7DB5056D5D75EABC7FFF5EAAAABEDF5257DAA8438EBA415568",
INIT_2A => X"4516D007FFFFFF1C042FB7D492A955C7F7FBD54380020ADA82BED57DF4508041",
INIT_2B => X"0870BAAA80070BAA2803DE00005F68A10BE802DB55E3DB555FFF68028ABA5D5B",
INIT_2C => X"00000000000000000000000000000125EFEBFFD2400EBFBFAFEFAA80070BAA2A",
INIT_2D => X"D53420BA082E82155AA802AAAAFF803DEBAAAFBC20BA55514000000000000000",
INIT_2E => X"5D04175EF0855575455D7BFFEAA5D5568ABAA2842AB55A28015545A284000BA5",
INIT_2F => X"FF7D57DE005D003DE00007FEAA10002ABFF450079C20BAAAAE9754500043DEBA",
INIT_30 => X"EFA2842AABA085768BFFA2AE820AAFF802ABEFAAFFEABEFAAFFFDEAA0051555E",
INIT_31 => X"E10F7D17FF5500000001008516AA10FFFFC01EF55556AB55F7D56AABAF7FBC01",
INIT_32 => X"75EFF7842AAAA5D7FD75EF087BFDFEF5D003DFEF002E95555F7FDD74BA08043D",
INIT_33 => X"EABFFAA84174BAAA80174AAAA86174AAAA843DE00087FE8A00F7843FF45AAFFD",
INIT_34 => X"0000000000000000000000000000000000000000000000001FFA2FFC2000A2FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000001000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"A1400802000020490000000000000240413C0A61590001D90213C90008510204",
INIT_02 => X"680108200010000054655C040080000041000000010402400800800009082011",
INIT_03 => X"00040100800020D0842240124210810043800504488000103081894288800000",
INIT_04 => X"00001410A00AA084000400C0060000040088323044201C850020820400101880",
INIT_05 => X"0200020040048A09202420000C00410402000025000800020804207000100800",
INIT_06 => X"10488704884D080202086A0A3429004012120004DC08125400A0008300821000",
INIT_07 => X"000800002C30204084381000128104000100002040003164040D800000400009",
INIT_08 => X"0440050003080202202400100080000000000C3E0408104C8000102300008810",
INIT_09 => X"4810240104111104200080120210A5104000A204615201500801010000AA10C0",
INIT_0A => X"81F525A82804010009029290200008B202238008080240000040100242048025",
INIT_0B => X"00A1141002C91844522A0004120488000800028000044000080020AF09240010",
INIT_0C => X"0408104081000810408100081040810008104040800408208040000008010121",
INIT_0D => X"4201E0B4000803200C150108008490809A002192462424202200440404204041",
INIT_0E => X"0804100160006000120002120499020A04A14650A32851962965190014200240",
INIT_0F => X"000000000080A200100021000000014020080021000000014020000014260082",
INIT_10 => X"0000000000000340080028000000014020080028000000014020008000008000",
INIT_11 => X"008000008000000000000081500010000100800000000000008C100080000012",
INIT_12 => X"05D0000880000006800058000020000000000005000000000000000048100100",
INIT_13 => X"0000D02E8040200000003401F80004000000000040026000274000900000001A",
INIT_14 => X"800023B8000030000000000042A00009AB00008800000000008012BA01001000",
INIT_15 => X"00A000106520350000040100000000000010C0200009BA000200000000000105",
INIT_16 => X"465196651B328CA8D26540544924272EB91004002022024048400000098030A0",
INIT_17 => X"6509425094250942509425094250942509425094250942509425094251946519",
INIT_18 => X"5094250942509425094250942519465194651946519465194651946519465194",
INIT_19 => X"2A05404808000000000000000014651946519465194651946519465094250942",
INIT_1A => X"69A69A69A68945B080201C92410480ABD102E689999E91BCD151200C30AE1C71",
INIT_1B => X"341A0D068341A0D068341A28A28A28A28A28A28A28A28A28A28A28A28A28A69A",
INIT_1C => X"FFC5B52068349A4D068341A0D269341A0D269341A0D068349A4D068349A4D068",
INIT_1D => X"0F7D17FFFFAAAE800000000000000000000000000000000000000000000003FF",
INIT_1E => X"EFAA843DE00F7803FEBAFFFFC2000557FEABEFA2D1400AA5D2AAAA00F7FFEAA1",
INIT_1F => X"4105555421EFF78028BEF5D003DFEFF7FFE8ABAF7802ABEFAAAE820000000021",
INIT_20 => X"AB45557BC0155007FFDEBAAA843DE00557BEAABAA2AEAABEFF78015555AA8017",
INIT_21 => X"154AAA2AA955FF00043DE005504175FF0851401455555555EFA2FBC01FFF7AAA",
INIT_22 => X"57DE105D2EBDF55557FFDE00552A974AAA2843DEAA5D2A820BA000428AAAAA84",
INIT_23 => X"517FFEFAAAEBDF45FFAEA8ABAF7D1400BAAAAE821EFF7D17DEAA5D2AAAAAA5D5",
INIT_24 => X"0000000000002ABFFA280154BAFF803DF45FFD17DFFFFFD56AA00557FC201000",
INIT_25 => X"4120ADA38E3F1EFA28F7DF7DFD7A2A4800000000000000000000000000000000",
INIT_26 => X"7A2A482038000A001C7A2803AE38FF843DEBAEBFFC20285D75EFBC7A2DB40082",
INIT_27 => X"C7EB8417555AA84104385D55421C7FF8028BEF41003FFD7F7F1EDA82F78E2DBD",
INIT_28 => X"5C7A2FBC51EFEBA0A8B6D5571C716D1475FFEAAA28E3FE385D71E8AAAAAA0A8B",
INIT_29 => X"50AA1C0428ABAB68E124BAA2AA955C708003FE285D00155FF0055451555D5F57",
INIT_2A => X"7FE825520ADA92495B7AE10412EBFF45497FFFE105D2E97482AA8038EAA412E8",
INIT_2B => X"F6DA284175C001000557FFEFB6A0BFF55F7AEAAA82FFDF40092B6A4871EFFFD5",
INIT_2C => X"0000000000000000000000000000028BEFA28E124AAF7843AF7DEBDB78FFFE3D",
INIT_2D => X"5517DF55A2FBC201008003DEAAA2D57FEAAF7FBFDF45AA800000000000000000",
INIT_2E => X"FFD57FE00FFAABFF45AA80020BA082E82155AA802AAAAFF803DEBAAAFBC20BA5",
INIT_2F => X"A5D5568ABAA2842AB55A28015545A284000BA5D5340145F78028BFF08003DF45",
INIT_30 => X"EF0855575455D7BD5555A2FBD75FFA2842ABFF5555575FF55557FEAAA2AABFEA",
INIT_31 => X"400A2802AABA002A954AA5D0028ABAF7AA820BAAAAE9754500043DEBA5D04175",
INIT_32 => X"2010FF80155EFF7D57DE005D003DE00007FEAA10002ABFF450079FFE005D2A97",
INIT_33 => X"2ABEFAAFFEABEFAAFFFDEAA00514200008517DFEFFF803FF45FFAAA8A00F7FBC",
INIT_34 => X"000000000000000000000000000000000000000000000028BFFA2AE820AAFF80",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000002000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033022000000180006",
INIT_01 => X"0000098218302849180060000C00424040000000080000080200090008510200",
INIT_02 => X"0801080200100000044008000080000041000000002002400800000009008010",
INIT_03 => X"0001000004000040000202000000000803006400088000003080040008C10000",
INIT_04 => X"0000100022008000000C08C00C00000400201830040000040000000400001820",
INIT_05 => X"0200000040000000248080210044000400000000000800000004000010000800",
INIT_06 => X"100007000049000202086A080000004010100000880800001000000030829000",
INIT_07 => X"000800002420000004201000128100000300002040003124040D802040400009",
INIT_08 => X"040005000108020220240020008000000000043E000000488000000100008811",
INIT_09 => X"0810040105111000202000024010A51040088080000000110000002000020084",
INIT_0A => X"040000000000010000040010200008B202230480080002000000100240008021",
INIT_0B => X"40003C020AC04400022808001000014000040088140000000000828000000820",
INIT_0C => X"0040004400044000040000400044000440000400002000221048840009012124",
INIT_0D => X"0002A00800000100440000000800800018002000008000800040022000000400",
INIT_0E => X"0804100100002000100002001001024800020001000080004000000800904000",
INIT_0F => X"000000000000A000102008000000014000082008000000014000000000240082",
INIT_10 => X"0000000000000240082001000000014000082001000000014000028000000000",
INIT_11 => X"028000000000000000000001400012000200000000000000000C100084000800",
INIT_12 => X"0000080000000004800000400020400000010000000000000000000048000000",
INIT_13 => X"0000900000010000000024080000000000000000000250002000200000000012",
INIT_14 => X"4000200000400000000000000290000100002000000000000000120000010000",
INIT_15 => X"0000001000000000010000000000000000104010000100000000000000000005",
INIT_16 => X"0000000001400080002100544924002A000004000020000080000000010032A0",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100400000000",
INIT_18 => X"0000000000000000000000000010040100401004010040100401004010040100",
INIT_19 => X"02A1410808000000000000000000000000000000000000000000000000000000",
INIT_1A => X"145145145146AB2A0CCC2A28A28A7AA0CDF0D1215281FC1A72E24C28E921AAA9",
INIT_1B => X"CA6532994CA6532994CA65145145145145145145145145145145145145145145",
INIT_1C => X"FFD9C63B95CA6532994CA6532B95CAE572994CA6532994CAE572B95CA6532994",
INIT_1D => X"FAAD1555FFF78400000000000000000000000000000000000000000000000200",
INIT_1E => X"AA5D2AAAA00F7FFEAA10F7D17FFFFAAAE801FF08557DF4555516AA00007BEABE",
INIT_1F => X"000557FC0010AAD57FF45A2D56AA0000043FFEFA2FFFDE1008556ABEFA2D1400",
INIT_20 => X"DEAA007FEAB45AAAE800AAF784020000000021EFAA843DE00F7803FEBAFFFFC2",
INIT_21 => X"421EFF78028BEF5D003DFEFF7FFE8ABAF7802ABEFAAAEA8BFF5D0415400F7FBF",
INIT_22 => X"015555AA80174105555401FF5D0415555557BFDFEF00517DE00A28028B450855",
INIT_23 => X"FFD7555AAD56AB45A2AE800AA5D7FFDEBAF7AEBDE00557BEAABAA2AEAABEFF78",
INIT_24 => X"000000000000155EFA2FBC01FFF7AAAAB45557BC0155007FFDEBAAA8417410AA",
INIT_25 => X"55556AA381C75EABEFBED1575C7E380000000000000000000000000000000000",
INIT_26 => X"81C516FBC7A2DB400824120ADA38E3F1EFA28F7DF7DFD7A2A4801EF085F7AF6D",
INIT_27 => X"38FF843DEBAEBFFC20285D75C0010AADF7AF6DB6D56FA3814003AFFFA2F1F8E3",
INIT_28 => X"BEF550412428F7F5FDE920875E8B45BEA0850BAE38002038000A001C7A2803AE",
INIT_29 => X"8E10AA802FB450851421C7FF8028BEF41003FFD7F7F1EDA82F78E2DBD7A2A4AD",
INIT_2A => X"E8AAAAAA0A8BC7EB8417555AA84104385D55401C75504125455575FAFD714557",
INIT_2B => X"5FFEAAA28E10438AAF5D2545BED56FB45BEA082082557BF8EBAF7AABFE385D71",
INIT_2C => X"00000000000000000000000000000175C7A2FBC51EFEBA0A8B6D5571C716D147",
INIT_2D => X"A80021FF007BE8BFF5D516AABA5D5568BEFF7D157555AA800000000000000000",
INIT_2E => X"5D002ABFFA2D16AAAA55517DF55A2FBC201008003DEAAA2D57FEAAF7FBFDF45A",
INIT_2F => X"A082E82155AA802AAAAFF803DEBAAAFBC20BA555140010AAFFE8BFFFFD17DEBA",
INIT_30 => X"00FFAABFF45AA803FFEF5500020BAFFD17DE10005568B55FF80154BAA280020B",
INIT_31 => X"1555D556AB555D5568A00AA843FF55085140145F78028BFF08003DF45FFD57FE",
INIT_32 => X"AAAAF7AABFEAA5D5568ABAA2842AB55A28015545A284000BA5D5342145550402",
INIT_33 => X"2ABFF5555575FF55557FEAAA2AA800AAAAD142155F7D57DF45FF8002010557FE",
INIT_34 => X"000000000000000000000000000000000000000000000015555A2FBD75FFA284",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000023FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B830084C1820E0000C36424840000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"000406A492E6E440842254D002108153422004800880000030C0315688C00006",
INIT_04 => X"00001201200090001205400000000094108C322644240C840008030440111800",
INIT_05 => X"222000444008010028404002A002009402400025080880000C04223000170900",
INIT_06 => X"12801628014B0B000A086CA6556800C012121004540816544522008200821100",
INIT_07 => X"1C08320054B624408428100094ADD080011721A04000316C140CA1A8A1F90019",
INIT_08 => X"00140500090B02C2E0EC04D1C08000000000647E858A104C920C81A5011088A6",
INIT_09 => X"40002481041F165820000101024061004004800567603592A801014C46426011",
INIT_0A => X"8404002020000101B0070310200008B60A23A51B28024CE24E40100260040004",
INIT_0B => X"2800340208811865D22BB384100E01090805A495100400050800E24D49A424C5",
INIT_0C => X"0C72A0872A0C72A0872A0C72A0C72A0872A0C595043950421400800009010104",
INIT_0D => X"4290A088812203360410110A400085539800210404C048CAC040464D28014405",
INIT_0E => X"0804101160006000101004A01811064B050204810240812241280D00200A0804",
INIT_0F => X"6D0141B0482A01AAEC3602330CD2A02952DC3502330CB4A0318B414000240082",
INIT_10 => X"5B4551630144C0155C3502330CD2A02952DC3602330CB4A0318B5600C587149B",
INIT_11 => X"FE04E587083B6A51005956308D1E8202C436375908AA840AD4513437640F1524",
INIT_12 => X"E020C67062F47B2872400044959BC42B1060F0D036B80B548523136C158878D8",
INIT_13 => X"8F0B27010A2699AAA3794392000D81852B0A050C224180062085134CD1719564",
INIT_14 => X"0AD57400C50500D94C8121713C02B555101C90705D71009604140C0418CE0C37",
INIT_15 => X"DC06A27C828E024D8C50965A40821568A06113801505010334AA73AA0666DAC2",
INIT_16 => X"04812048123408C0822040004C248604B2100400100084008001D0113920060C",
INIT_17 => X"4812048120481204812048120481204812048120481204812048120481204812",
INIT_18 => X"8020080200802008020080200812048120481204812048120481204812048120",
INIT_19 => X"00A0014200000000000000000020080200802008020080200802008020080200",
INIT_1A => X"4104104104140D220A4A380000002A80E900C4C1100830181621409C80210821",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000410",
INIT_1C => X"FFC1F83800000000000008040000000000000000000201000000000000000000",
INIT_1D => X"0F7842AA00002A80000000000000000000000000000000000000000000000200",
INIT_1E => X"4555516AA00007BEABEFAAD1555FFF784020AAF7D542155F7D1400AAF7FFFDE0",
INIT_1F => X"FFFAAAEA8ABAFFD17FEBAFFAA800AA007FFDFFFA28428A000000001FF08557DF",
INIT_20 => X"00AAF78028AAAFF84020AAFFFBEABEFA2D1400AA5D2AAAA00F7FFEAA10F7D17F",
INIT_21 => X"40010AAD57FF45A2D56AA0000043FFEFA2FFFDE1008556AB45555568A10A2FFC",
INIT_22 => X"03FEBAFFFFC2000557FC0155FFD1555FF0804000AA000428A10AAAA801EFFFD1",
INIT_23 => X"8428A10087FD7400552EBDFEFA2FBFFF550000020000000021EFAA843DE00F78",
INIT_24 => X"00000000000028BFF5D0415400F7FBFDEAA007FEAB45AAAE800AAF78428B45A2",
INIT_25 => X"E3DF450AAF7F1FDE38FF8A2DA101C2A800000000000000000000000000000000",
INIT_26 => X"01C0E001EF085F7AF6D55556AA381C75EABEFBED1575C7E380000BAF7DB4016D",
INIT_27 => X"38E3F1EFA28F7DF7DFD7A2A4AFABAFFDF7AE82F7AA870AA0071F8FFFBE842DA1",
INIT_28 => X"B455D5B68A28A2FFC20AAEB842DAAAE38A02082E3FBEFBC7A2DB400824120ADA",
INIT_29 => X"8A28AAA4801FFE3DF40010AADF7AF6DB6D56FA3814003AFFFA2F1F8E381C516D",
INIT_2A => X"001C7A2803AE38FF843DEBAEBFFC20285D75C2145F7DF525EF140A050AA1C002",
INIT_2B => X"0850BAE3802DB6DAA8A28A00007FD74284120BFFFFBEF1F8F7D080A02038000A",
INIT_2C => X"000000000000000000000000000002DBEF550412428F7F5FDE920875E8B45BEA",
INIT_2D => X"A80020BAFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE10552E8000000000000000",
INIT_2E => X"085568BEFF7803FE10552E821FF007BE8BFF5D516AABA5D5568BEFF7D157555A",
INIT_2F => X"5A2FBC201008003DEAAA2D57FEAAF7FBFDF45AA803FEBAFFFBEAA00F7AE974BA",
INIT_30 => X"FFA2D16AAAA55517DF55557FEAAAAA2FFC00AAAA803FEAAA2AA82000A2FFFDF5",
INIT_31 => X"1EF552E974BA550028ABAA280001FFAAFFC0010AAFFE8BFFFFD17DEBA5D002AB",
INIT_32 => X"ABFF082E820BA082E82155AA802AAAAFF803DEBAAAFBC20BA555142155F7FFC0",
INIT_33 => X"7DE10005568B55FF80154BAA2803FFFFA2AAAAA00007FD74BA08003DFFFFFD16",
INIT_34 => X"00000000000000000000000000000000000000000000003FFEF5500020BAFFD1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000002000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C048000C048400380000007026040000000080000088200002802153231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"210D050012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"0080100022408000060DE0000066630C70241827041000040800820480001AA4",
INIT_05 => X"0240000C400000003C808003E0C8001401000000040900020904004000070800",
INIT_06 => X"1800068000491300CF0969A421C0004018184000100804005784000130821200",
INIT_07 => X"7E8C53200CA4850224301807D1CB45900147E03040083124FC0CD0C8A1FF0019",
INIT_08 => X"0046050013081206A4A503A9E8C0812000001C7E11A24058B84D40E33992D98F",
INIT_09 => X"010004810491175C20000080000821004010C01086003C13E000004EDF020400",
INIT_0A => X"000000000000010000180018200408B27E234913E9000CFA09A8180248001000",
INIT_0B => X"ACA0141000800021826933E03662802B3001E09F000000023000000000000867",
INIT_0C => X"0832F0C32F0832F0832F0C32F0832F0832F0C197861978400000000208010100",
INIT_0D => X"05FA0201E7F3F01F40401C17E800C7F3380020000000006AE01180493C5BC1AF",
INIT_0E => X"000200F500002200004005002001408400000000000000000000053A4096F807",
INIT_0F => X"246FC1B17B2C53F2FC16691DB587201EDDF4162B1DB527201EDDC46070241001",
INIT_10 => X"2A67DF2A01D5CC9794162B1DB587201EDDF416691DB527201EDDD884272592D6",
INIT_11 => X"288007258E995D5A825DBA569F9FF02547068618CD3CC45B7863AE7EC00D4B12",
INIT_12 => X"F6208C6CCA5C33717461C045B5B182019473D19D7CCD856106F31A683621BDFC",
INIT_13 => X"866E2FB10A652CC8E3538BBA01624E51AA6C0469AC5493F5688532966471A9C5",
INIT_14 => X"4F9B740041E1F5759001B4AA1853E6D5144AA9C914C8608D2724A4C4118D992B",
INIT_15 => X"DE07EAD9825682D4A36C0B0B4B85112B2C4A05D3E6D5051893335EB0072AA85A",
INIT_16 => X"00000000008000000821000048260020000004001DC0800000010E7F70171401",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0100401004010040100401004000000000000000000000000000000000000000",
INIT_19 => X"2A21010808000000000000000000401004010040100401004010040100401004",
INIT_1A => X"4924924924890380800016A28A28802B10B83728C1111026C152A23010848658",
INIT_1B => X"6432190C86432190C86432082082082082082082082082082082082082082492",
INIT_1C => X"FFDE003AC964B2592C964B2592C964B2592C964B2592C964B2592C964B2592C9",
INIT_1D => X"5FFAA80155F78400000000000000000000000000000000000000000000000200",
INIT_1E => X"55F7D1400AAF7FFFDE00F7842AA00002AAAA10FF8002155F7FFC200008041755",
INIT_1F => X"5FFF7842AB55080000145557FE8AAA080000155F7FFFDEAA0000020AAF7D5421",
INIT_20 => X"2000FF80020AAA2AAAABFF002E801FF08557DF4555516AA00007BEABEFAAD155",
INIT_21 => X"A8ABAFFD17FEBAFFAA800AA007FFDFFFA28428A00000028B4555043DFFFFFAE8",
INIT_22 => X"FEAA10F7D17FFFFAAAE80000A284174AAFF8428AAAFF8415545AAFBD7545F7AA",
INIT_23 => X"00000105D55400AA082A82155F7FFFDEAA08556ABEFA2D1400AA5D2AAAA00F7F",
INIT_24 => X"0000000000002AB45555568A10A2FFC00AAF78028AAAFF84020AAFFFBC215508",
INIT_25 => X"E3F5C000014041256DEBA487145F784000000000000000000000000000000000",
INIT_26 => X"2080E000BAF7DB4016DE3DF450AAF7F1FDE38FF8A2DA101C2AAFA00EB8E0516D",
INIT_27 => X"381C75EABEFBED1575C7E3802FB551C0E0516D417FEDA921C000017DEBF5FDE9",
INIT_28 => X"B55410A3FFC7F7A087000FF80070BAAAAAADBD70820801EF085F7AF6D55556AA",
INIT_29 => X"556DA2FBD7545F7AAAFABAFFDF7AE82F7AA870AA0071F8FFFBE842DA101C0E2D",
INIT_2A => X"400824120ADA38E3F1EFA28F7DF7DFD7A2A480000BE8A17482F78A28A92E3841",
INIT_2B => X"A02082E3FBC217D1C0E0500041554508208208017DF7F5FDE9208556FBC7A2DB",
INIT_2C => X"000000000000000000000000000002DB455D5B68A28A2FFC20AAEB842DAAAE38",
INIT_2D => X"52EBDE00AAAE975FFAAD1420005504001FFAA8015545F7800000000000000000",
INIT_2E => X"5504001FFAAD17DE00082E820BAFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE105",
INIT_2F => X"F007BE8BFF5D516AABA5D5568BEFF7D157555AA803DF45552E975EF007FFFE00",
INIT_30 => X"EFF7803FE10552EBDF45002EBFF55FF8017410FF84154BAAAAABFF450000021F",
INIT_31 => X"400F7AEA8A10A284175FFAAFBD5555F7AEBFEBAFFFBEAA00F7AE974BA085568B",
INIT_32 => X"DE1008517DF55A2FBC201008003DEAAA2D57FEAAF7FBFDF45AA8002000FFAE95",
INIT_33 => X"C00AAAA803FEAAA2AA82000A2FFC21EF552A954100851554000004021FFFFD17",
INIT_34 => X"00000000000000000000000000000000000000000000003DF55557FEAAAAA2FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00010100926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"0004122122029100100C00001200009C40A83A2044360C84190BAC04E0101820",
INIT_05 => X"027000004009050064C8C00104C10184034010250089C00EB004327064B60900",
INIT_06 => X"1B9416B94149000402086D42142800C012125804440812541027008230821380",
INIT_07 => X"0008320014B02848A4A8100015C55500057801A04000712C040CB1F880600009",
INIT_08 => X"005005000908020220E40170008042000000557E048A144C800590010000882D",
INIT_09 => X"0100250104B5310020000100020821004016CC1C616401910801010100CA2040",
INIT_0A => X"800000000000010192072310200028B6022346080802C0074AC0100259001004",
INIT_0B => X"A8201410008088C5D2288004120E802908800488000500050800404D49A42EB0",
INIT_0C => X"0400000000040000000000000040000000000000020000000000000008010102",
INIT_0D => X"4A02008000000360401021280800E400B800610C844848200028448400000000",
INIT_0E => X"000000086000600040D045E4195104D5854284A14250A12A512A880828984008",
INIT_0F => X"85D480949E07A80948354B6E68982167061037496E6838216706206810240000",
INIT_10 => X"652138E510B456587037496E689821670610354B6E6838216706220431961CA9",
INIT_11 => X"C2043196186A91674011CE61403562274AA49CD594CF00039C7C414B6509DA22",
INIT_12 => X"8A2E6A983014780CC8604040424A5323845932E620295879818170304B2F5002",
INIT_13 => X"8F019451654B9104A328665603148895D44E0251142B42A3D8B2A5C882519432",
INIT_14 => X"0AC5DC06A6C6A465AA0091482382B17614F2202858EE300991415B45CD530602",
INIT_15 => X"4000052E08DC8047F17D1C7C3C02128E587D6A02B17605A130A4E8BF00225885",
INIT_16 => X"84A1284A123508508220808048240604B2100C00022084809000D000393722A1",
INIT_17 => X"4A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A12",
INIT_18 => X"A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A128",
INIT_19 => X"F1228154000000000000000000284A1284A1284A1284A1284A1284A1284A1284",
INIT_1A => X"75D75D75D75FFAFEFEFEEEAAAAAAFBF3FC1FF77DDFE7EFBEFFE7CFC0044FBEFB",
INIT_1B => X"FAFD7EBF5FAFD7EBF5FAFD75D75D75D75D75D75D75D75D75D75D75D75D75D75D",
INIT_1C => X"FFC0003BF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5",
INIT_1D => X"F007FE8A00AAFBC0000000000000000000000000000000000000000000000200",
INIT_1E => X"55F7FFC2000080417555FFAA80155F7842AB55552E821FFFFD5555EF552ABDFE",
INIT_1F => X"A00002A821EF5D7BC21FFFFFBD55EFAAD1554BA00556AA00AAD16AA10FF80021",
INIT_20 => X"FF45A2AABFEBA082A975555D55420AAF7D542155F7D1400AAF7FFFDE00F7842A",
INIT_21 => X"EAB55080000145557FE8AAA080000155F7FFFDEAA00002AB45082A821EF5D557",
INIT_22 => X"BEABEFAAD1555FFF7842AABAA2FFE8BEF5D517FF455D554214500043DEBAAAFF",
INIT_23 => X"AABDF555D2E955EFA28428A10552EBFEAAAAD1401FF08557DF4555516AA00007",
INIT_24 => X"00000000000028B4555043DFFFFFAE82000FF80020AAA2AAAABFF002E80000AA",
INIT_25 => X"EBD5525C74124B8FC71C71EFA28AAF5C00000000000000000000000000000000",
INIT_26 => X"8AAD16FA00EB8E0516DE3F5C000014041256DEBA487145F78428B6D4120851FF",
INIT_27 => X"AAF7F1FDE38FF8A2DA101C2A871C74975C01FFEBF5D25EFA2D555482085F6FA2",
INIT_28 => X"B7D1C24851FF495F7FF55A2A0BFE921C2E9557D415B400BAF7DB4016DE3DF450",
INIT_29 => X"214508003FEAABEFFEFB551C0E0516D417FEDA921C000017DEBF5FDE92080E2A",
INIT_2A => X"7AF6D55556AA381C75EABEFBED1575C7E38028A82B6F1E8BFF495F78F7D49554",
INIT_2B => X"AADBD7082087000AAA4BFF7D5D20905C7AA842DA00492EBFEAABED1401EF085F",
INIT_2C => X"000000000000000000000000000002DB55410A3FFC7F7A087000FF80070BAAAA",
INIT_2D => X"78028BFF0004175EFA2D54214508042AB455D517DEBAA2D54000000000000000",
INIT_2E => X"AAD557410007BFDEAAA2D57DE00AAAE975FFAAD1420005504001FFAA8015545F",
INIT_2F => X"AFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE10552E975450051401EFA2D5421EF",
INIT_30 => X"FFAAD17DE00082EA8BFF5504175FF087BFFF45AA843FE005D2A955FF087BC20B",
INIT_31 => X"BFF087BEABEF00554215500003FEBAFFFBFDF45552E975EF007FFFE005504001",
INIT_32 => X"FEAAFFD5421FF007BE8BFF5D516AABA5D5568BEFF7D157555AA8028A00FFD16A",
INIT_33 => X"17410FF84154BAAAAABFF45000017410AA803DFEF550402155A2843FE00082AB",
INIT_34 => X"00000000000000000000000000000000000000000000003DF45002EBFF55FF80",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000033FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"000103A7A00904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000120122009000100C00000000000400A83A2044200C840000800400101820",
INIT_05 => X"020000004008010024C0C0010040000402000025000800020004207000100800",
INIT_06 => X"108016080149080002086807542800C012120004440812541020008230821000",
INIT_07 => X"4008120054B42850B42A100010ED1500010001A040003164040CF5E201400009",
INIT_08 => X"00400500090A020220A40A7000800000000014FE8508144C924080C100008801",
INIT_09 => X"0000040104111100200001000200210040008004616001910801010000422000",
INIT_0A => X"800000000000010190070310200008B202236D080802400002C0100240000000",
INIT_0B => X"0000141000800844522800041204000008000488000400000800004D49240820",
INIT_0C => X"0400004000000000000004000000000000004000000000000000000008010100",
INIT_0D => X"42020080000002204010010808008000B8002104044048200000440400000000",
INIT_0E => X"0000000000006000000000201811004005020481024081224128080820984000",
INIT_0F => X"CBA340480040A100A42008000161C140000420080001C1C14000032010240000",
INIT_10 => X"1A8A039600022260042001000161C140000420010001C1C140001604E8084341",
INIT_11 => X"1E04E8082580E2B8802201014800C220A21829A302F1C024010C001124020C8C",
INIT_12 => X"0024ACA60CA000048228404401004418012787124648157780120B8678C00080",
INIT_13 => X"00009001072D04730000241000CB1325E78E0186030240000083B60239800012",
INIT_14 => X"00001001EF6F4163C480481506800004000CFD55196CB012481812049495C194",
INIT_15 => X"40068248800108B8FB61A0401200845594965000000400568D0CFB7800550605",
INIT_16 => X"04812048123408408220000048240604B210040000008400800B0000090022A1",
INIT_17 => X"4812048120481204812048120481204812048120481204812048120481204812",
INIT_18 => X"8120481204812048120481204812048120481204812048120481204812048120",
INIT_19 => X"2820014000000000000000000020481204812048120481204812048120481204",
INIT_1A => X"3CF3CF3CF3CFFBBEEEEEFE79E79EFAABDDFAF369CB91FE1EF7D3AEBBDBAFBEFB",
INIT_1B => X"FE7F3F9FCFE7F3F9FCFE7F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"FFDFFFC1FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"AAAAEAAB45082E80000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFD5555EF552ABDFEF007FE8A00AAFBE8BEFA2D568ABA00003DF555555574A",
INIT_1F => X"155F78428AAA007FE8A1008002AABA555155400557BC2010557BEAB55552E821",
INIT_20 => X"FFFF082EBDEBAA2D1420105D002AA10FF8002155F7FFC2000080417555FFAA80",
INIT_21 => X"C21EF5D7BC21FFFFFBD55EFAAD1554BA00556AA00AAD140145AA8028ABA002EB",
INIT_22 => X"FFDE00F7842AA00002A80155A2AEA8A10080428A10FFAEBFFEF5D0428B45A2FF",
INIT_23 => X"5568A000000175FFF7D155545F7FBC0010FFAA820AAF7D542155F7D1400AAF7F",
INIT_24 => X"0000000000002AB45082A821EF5D557FF45A2AABFEBA082A975555D55400BA00",
INIT_25 => X"000E38F6D4155504AAA2AEAAB6D0024800000000000000000000000000000000",
INIT_26 => X"05D75E8B6D4120851FFEBD5525C74124B8FC71C71EFA28AAF5E8BFFB6D56DA82",
INIT_27 => X"0014041256DEBA487145F78428ABA147FEDA10080E2AAAA555552400417FC200",
INIT_28 => X"155BE8028A82002EB8FC70024BAEAAB6DB4202849042FA00EB8E0516DE3F5C00",
INIT_29 => X"DFD7550428B55A2F1C71C74975C01FFEBF5D25EFA2D555482085F6FA28AAD147",
INIT_2A => X"4016DE3DF450AAF7F1FDE38FF8A2DA101C2A80145B6AEA8A10080E2DA00F7A0B",
INIT_2B => X"E9557D415B400AA00556DA000004175FFE3D15757DE3F5C0038FFAA800BAF7DB",
INIT_2C => X"000000000000000000000000000002AB7D1C24851FF495F7FF55A2A0BFE921C2",
INIT_2D => X"2D568BEFFFD57FE10002AAABEF0051400AAA2AAAABFF08000000000000000000",
INIT_2E => X"5D5142000007BC20105D5568BFF0004175EFA2D54214508042AB455D517DEBAA",
INIT_2F => X"0AAAE975FFAAD1420005504001FFAA8015545F78028AAA557FFFE00082EAAAAA",
INIT_30 => X"10007BFDEAAA2D557555FF8028A00082EAAB45000028ABAFFFBC20AA08043DE0",
INIT_31 => X"A10002ABFE00F7803FF555D002AB55AAD1575450051401EFA2D5421EFAAD5574",
INIT_32 => X"20BAFFAE820BAFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE10552E82155FFAAA8",
INIT_33 => X"FFF45AA843FE005D2A955FF087BC20AA00517DE000804175EFAAD1555EFA2D14",
INIT_34 => X"000000000000000000000000000000000000000000000028BFF5504175FF087B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000080000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"0001100024A0800000440000000000040088322044200C840000011400151800",
INIT_05 => X"A200014C4000000020000000000B8094020000254C8800000514203000108800",
INIT_06 => X"10000600004B0044020868021428004012120005540812540020008600831000",
INIT_07 => X"00086100043224489428100010811100010001A040003124040CAC6000400009",
INIT_08 => X"00160500090A0282A06400100080C300000005BE0488104C8000000100008800",
INIT_09 => X"00000581041110022000000002002100400080046140011008010100008A0400",
INIT_0A => X"800000000000010180060210200008B2022304080800400007C0100240000000",
INIT_0B => X"0004140000800844522800041004000008000080000400000800000D09240000",
INIT_0C => X"0400004000040000400000000000000000004000020000200000000008010100",
INIT_0D => X"4A00008000000260001001280000C400B0002000000000000000440400000000",
INIT_0E => X"0000000840006000000000001001004004000000000000020100000000000000",
INIT_0F => X"0000000000000000002021000000000000002021000000000000046000240000",
INIT_10 => X"0000000000000000002028000000000000002028000000000000020000008000",
INIT_11 => X"0200000080000000000000000000020001008000000000000000000004000012",
INIT_12 => X"0020000880000000006000400080C0000000000D081202800000000000000000",
INIT_13 => X"0000000100402000000000100000040200100000000000000080009000000000",
INIT_14 => X"0000100000003088014000000000000400000088221100000000000401001000",
INIT_15 => X"4000000800000000048407170500000000000000000400000200000000000000",
INIT_16 => X"00000000023000000220000048240404A010040000008000000000000000020C",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0020014000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000020000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFC0000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"555003DE10A2FBC0000000000000000000000000000000000000000000000200",
INIT_1E => X"BA00003DF555555574AAAAAEAAB45082EBFE000004020AA552E80000F7FBC214",
INIT_1F => X"A00AAFBFDEBA555568BEFA2FBE8A10F7802AA0055003FE10007BE8BEFA2D568A",
INIT_20 => X"55EFF78428BEFAAD17DF55AAAEAAB55552E821FFFFD5555EF552ABDFEF007FE8",
INIT_21 => X"28AAA007FE8A1008002AABA555155400557BC2010557BFFFEFA2FFC20005D2A9",
INIT_22 => X"417555FFAA80155F7843DF455D2AA8B45AAD57FF55A2FBC21FFA28415400FF80",
INIT_23 => X"514200055002AA00AA802AABA002E9740055516AA10FF8002155F7FFC2000080",
INIT_24 => X"00000000000000145AA8028ABA002EBFFFF082EBDEBAA2D1420105D003FFFF08",
INIT_25 => X"412A87010E3F5C0145410E3DE28B6FFC00000000000000000000000000000000",
INIT_26 => X"8147FE8BFFB6D56DA82000E38F6D4155504AAA2AEAAB6D0024B8E381C0A00092",
INIT_27 => X"C74124B8FC71C71EFA28AAF5F8EAA495F68BFFA2F1EFA38E38428A005D0038E2",
INIT_28 => X"FFFBEF5C0000492A955FFF78428BEFB6DB7DF45AAAEA8B6D4120851FFEBD5525",
INIT_29 => X"21EFAA8E10400E38E28ABA147FEDA10080E2AAAA555552400417FC20005D75F8",
INIT_2A => X"0516DE3F5C000014041256DEBA487145F7843FF7D4120A8B6DAAD17FF55B6F5C",
INIT_2B => X"B4202849043FFC7005F4501041002FA38A2842AA82142095428415F6FA00EB8E",
INIT_2C => X"0000000000000000000000000000007155BE8028A82002EB8FC70024BAEAAB6D",
INIT_2D => X"8002AAAA5D2A82000082E95400A2D542155002ABDEBAF7FBC000000000000000",
INIT_2E => X"A2802AA105D002AABA5D7BE8BEFFFD57FE10002AAABEF0051400AAA2AAAABFF0",
INIT_2F => X"F0004175EFA2D54214508042AB455D517DEBAA2D56AABA087BEABEFAAD57DEAA",
INIT_30 => X"00007BC20105D556ABFFF7D142010082A955EFFF8428BFFFFFBFDF55A2AEA8BF",
INIT_31 => X"BEFA2D57DF45F7D1401FFA2AA82000AAAAA8AAA557FFFE00082EAAAAA5D51420",
INIT_32 => X"54AA007BFDE00AAAE975FFAAD1420005504001FFAA8015545F7803FFEF08002A",
INIT_33 => X"AAB45000028ABAFFFBC20AA08043FF55087BD740000043DEAAA2842AA005D001",
INIT_34 => X"000000000000000000000000000000000000000000000017555FF8028A00082E",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000003000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"010108A802BB00080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"8BFA58800005C40A46240252145148B38248030356415A4E62B6FC660F287240",
INIT_05 => X"0F05EA11E570000D610000000710296E542B6E3A825C15FB30A643695BFC2D56",
INIT_06 => X"00000200021100C87570B08224C8AB52C0A8030140BCC0460050690A95C8383D",
INIT_07 => X"76F500240510A00205F0A407D0021A155378900002A002433A0AA00EE6E79564",
INIT_08 => X"00015995440C8327241440096A2800002828123D542910380004E03103624040",
INIT_09 => X"0010222D90409A05B2CB2CA400200209E5601044A24000000462A60018880100",
INIT_0A => X"300000000000259200140001A15000017F0051D0F837248C005514AC40C08205",
INIT_0B => X"395012004240014891801000495D40192D100000000005452D54000C09070003",
INIT_0C => X"6110001100011000110001100011000110001080008800080005202280801080",
INIT_0D => X"BB4000140A80A5C8000102ED0044008004AD324000000008003561180063DB4F",
INIT_0E => X"1400404912AA28AA890BA00000024800480000000000000200802151025062C0",
INIT_0F => X"6D0031F554E11C596A64003195933741477264003195555B418687E358360208",
INIT_10 => X"41CD50A499CF47DCB264003195933741597264003195555B4198843940076D29",
INIT_11 => X"043D400758486A556489347FE5F409CBC1362510695B6288743123C952518520",
INIT_12 => X"B1C74424EAE2992046EB70026486035600CEC45CBCA809654B48163CCC895E1E",
INIT_13 => X"C383298E3A242DEA151848302BFD6D522B10C7EC71F6C1DB071D1216E078C4C1",
INIT_14 => X"8B93D037DAAABC982BE22267A2E2E4F44AA1DC5E37400C9EE1B7B638E8849D23",
INIT_15 => X"86E6A2EE015998B28654565A003F0068E35352C1CAE48BFBF3A6C9B7B286B4DA",
INIT_16 => X"00000000009000040A8000452110A8442040D655602A102A0027E2C423202840",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"B020000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"28A28A28A28F4EF2FC3C34F3CF3C2AC31DF7A22A898D21B4C9838D30B6A7B451",
INIT_1B => X"F4FA3D3E8F4FA3D3E8F4FA68A68A68A68A68A68A68A68A68A68A68A68A68A28A",
INIT_1C => X"FFC00003E9F4FA7D3E9F47A3D1E8F47A3D1E8F47A3D3E9F4FA7D3E9F4FA7D3E9",
INIT_1D => X"AFF80001FF002A80000000000000000000000000000000000000000000000200",
INIT_1E => X"AA552E80000F7FBC214555003DE10A2FBC21FFFFFBFDF45A2D56AB45FFFFD54B",
INIT_1F => X"B45082E974BA5D7BFDF55A2FFFFE005D7BC0010002E954AA087FFFE000004020",
INIT_20 => X"7410FFD1555550000020BAAAFFE8BEFA2D568ABA00003DF555555574AAAAAEAA",
INIT_21 => X"BDEBA555568BEFA2FBE8A10F7802AA0055003FE10007BC0000082A9740055001",
INIT_22 => X"ABDFEF007FE8A00AAFBD55EFAAFBD74105504021FF5D2EAAABAFFFBD55FF002A",
INIT_23 => X"517DF45AAFFFFEAAFFAABFE10007FC00AA087FEAB55552E821FFFFD5555EF552",
INIT_24 => X"0000000000003FFEFA2FFC20005D2A955EFF78428BEFAAD17DF55AAAE820AA5D",
INIT_25 => X"AADB6FB6DFFFBD54AAE38E021FF0824800000000000000000000000000000000",
INIT_26 => X"A1C7FF8E381C0A00092412A87010E3F5C0145410E3DE28B6FFC21C7E3F1F8F55",
INIT_27 => X"6D4155504AAA2AEAAB6D002492482497BFDF45AAFFF8E385D7BC5000002E904B",
INIT_28 => X"010142E90428490015400FFDB555450804070BABEF5E8BFFB6D56DA82000E38F",
INIT_29 => X"DAAAFFF1D55FF002EB8EAA495F68BFFA2F1EFA38E38428A005D0038E28147FC2",
INIT_2A => X"851FFEBD5525C74124B8FC71C71EFA28AAF5D25D7B6F1D54384904021FF5D2AA",
INIT_2B => X"B7DF45AAAE820925D5B7DF45A2F1FDEAAEBAABDE001471C20921475E8B6D4120",
INIT_2C => X"0000000000000000000000000000038FFFBEF5C0000492A955FFF78428BEFB6D",
INIT_2D => X"7FBC2145AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF00000000000000000000",
INIT_2E => X"557FD7410082A800AA557BEAAAA5D2A82000082E95400A2D542155002ABDEBAF",
INIT_2F => X"FFFD57FE10002AAABEF0051400AAA2AAAABFF080000000087BFDF55A2FFE8AAA",
INIT_30 => X"105D002AABA5D7BC20005D2E800BA080417400F7FBD75450800174AAFFD168BE",
INIT_31 => X"4AA0800001EF5D2ABDEBAF7D1575EF082EAAABA087BEABEFAAD57DEAAA2802AA",
INIT_32 => X"0000555568BFF0004175EFA2D54214508042AB455D517DEBAA2D540155F7D155",
INIT_33 => X"955EFFF8428BFFFFFBFDF55A2AE82010557FFDF55A2D57FEAAAAAEBFE1055514",
INIT_34 => X"00000000000000000000000000000000000000000000002ABFFF7D142010082A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000001000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"294ADB4AFFCBF0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"DB7A40806FE4040840EBC563A0150A0926146FECB04196482236FC2005282AE1",
INIT_05 => X"0403DA0383200831C68206D7E6D0250834336D1E81500FDB306045255BFC2076",
INIT_06 => X"D0002200022D1C59E53558D3EBFC6701CBC303163670497AFF00291B3C0E2015",
INIT_07 => X"F81684248A38B022475DCA9BD00116E33CC3821774BB55F53BB42329AA3C0CEA",
INIT_08 => X"1660700CE0641527241060AD844E1C0088001223022D189A2800542219204903",
INIT_09 => X"B6D94C1C1C51DFF881861CBE0305A12A0321810217C01D34EDC98FFA1C8E0000",
INIT_0A => X"F1F1FD8F8FBDE40E001E000B3A5DAADAFDDA5DA79350DF70027CE86F047BEF19",
INIT_0B => X"2DD8141817C00319F8E853E64D73A08BFF00E9A7415606747E6610052CDEE97F",
INIT_0C => X"4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A7800617112E46F05D0",
INIT_0D => X"BFF252D4CFEB69FF7A5F5AFFCCA787F7FE67C2180000006CE8A3F06ABD73DBCF",
INIT_0E => X"94BB02C9F99FD0678B87A0003000D8D02E00000000000000040025D3C21463D6",
INIT_0F => X"6D2BF232221ABD9CA854DFDD64A67D42C0F054DFDD64667D42C063E57A8F7B45",
INIT_10 => X"EFBB5AEDAA504801F054DFDD64A67D42C0F054DFDD64667D42C07237DFE5865F",
INIT_11 => X"3A33DFE58EAE7F5AB50D0806A9A2E0DFFF47DEDC496DA3181A0CC71440F9FBC3",
INIT_12 => X"7056E9C9C3FC95949AEFF556EF9C75E7DCF1EB1B6E6FCDC87CB35FC94B36AECF",
INIT_13 => X"92B29382AF5B6AAAE594A4C0DBFDAD94AA669809809FEFAF4157ADB55572CA52",
INIT_14 => X"BEBF41AE33F32ADD543430808BABAF50E1A5EB4BAEA45A250202FE0ADD39387F",
INIT_15 => X"E83FB669523E865D4B1293AB6B90BF2F0E30EDEFAFD0B3FBD72E9E90D20A003F",
INIT_16 => X"0000000002F840000BCE0B6F67B3F845E017C833F6AAC02B002A2EFF22D4073D",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"CC0C006000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"34D34D34D352324C3434C0EBAEBA21BBE5F04006013DB9880A5D25C3230B88A7",
INIT_1B => X"1A0D06A351A0D06A351A0D34D75D34D34D75D34D75D34D34D75D34D75D34D34D",
INIT_1C => X"FFC00002351A8D46A351A8D46A351A8D46A351A8D468341A0D068341A0D06834",
INIT_1D => X"0007BEAB55FFAA800000000000000000000000000000000000000000000003FF",
INIT_1E => X"45A2D56AB45FFFFD54BAFF80001FF002A821FFFFFFFFFFFFFFBFDFEFAAD14201",
INIT_1F => X"E10A2FBEAB45A28000010082A975EFA2D140145007BC21FF5D2A821FFFFFBFDF",
INIT_20 => X"54AA0855575FFAAD57FE005D7BFFE000004020AA552E80000F7FBC214555003D",
INIT_21 => X"974BA5D7BFDF55A2FFFFE005D7BC0010002E954AA087FD7400082E954AA08001",
INIT_22 => X"5574AAAAAEAAB45082EBFFFFF7D16AB45FFFFEABEF007BD74005555555EFF7AE",
INIT_23 => X"84154BA082E801FFAAFBC0155555568B45552EA8BEFA2D568ABA00003DF55555",
INIT_24 => X"00000000000000000082A97400550017410FFD1555550000020BAAAFFC0145AA",
INIT_25 => X"F7F1FAFD7A2D5400001C7BEDB7DEBA4800000000000000000000000000000000",
INIT_26 => X"F4124821C7E3F1F8F55AADB6FB6DFFFBD54AAE38E021FF0824851FFFFFFFFFEF",
INIT_27 => X"10E3F5C0145410E3DE28B6FFEFB45AA8E070281C20925FFBEDB451451C7BC01E",
INIT_28 => X"4280024924AA1404174AA0055505EFBEDB7AE385D7FF8E381C0A00092412A870",
INIT_29 => X"54005D5B575EFEBAE92482497BFDF45AAFFF8E385D7BC5000002E904BA1C7FD5",
INIT_2A => X"6DA82000E38F6D4155504AAA2AEAAB6D0024BFFD7FFDB6AB7DFFF5EDBC71C7BD",
INIT_2B => X"4070BABEF5C516DAA8A124921C20801FFB6F5C0145555B68B7D4124A8BFFB6D5",
INIT_2C => X"0000000000000000000000000000002010142E90428490015400FFDB55545080",
INIT_2D => X"000155FFF7FBFDFEFFFD568B45AAD5400005D7BFFFEFAA800000000000000000",
INIT_2E => X"FFFFD5545557BC21FF080002145AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF0",
INIT_2F => X"A5D2A82000082E95400A2D542155002ABDEBAF7FBFDF55A2AA974AA5D04001EF",
INIT_30 => X"10082A800AA557BD74BA0004000AA5500174AA0855421FFFFFBEAAAA5D7BEAAA",
INIT_31 => X"BFFF7D57FF455D7FD54105D7BD75FFAAAA80000087BFDF55A2FFE8AAA557FD74",
INIT_32 => X"8BEF000028BEFFFD57FE10002AAABEF0051400AAA2AAAABFF08003FF55F7FFEA",
INIT_33 => X"17400F7FBD75450800174AAFFD1555FFA2AA800105504001EFFFD140145557BE",
INIT_34 => X"0000000000000000000000000000000000000000000000020005D2E800BA0804",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000033FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"0405D434003F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"50805AC31007D6125724029216554A9847669903D640EC8E2001002604503004",
INIT_05 => X"07008000E0EA11803850C800010022660C1C0065003C0404002646DC20A02D40",
INIT_06 => X"30A03A0A138900001127A09234C81FF040000000002C44D620F0228454C83810",
INIT_07 => X"405584280B10014003A8067400920810FF3C72024300A0030048221ACEE383E4",
INIT_08 => X"1000C983E6041505253500F66E620428000B1804000152E52801A20200840900",
INIT_09 => X"0820500B90419005B0C309402030060860E01004A828408800440405E3502940",
INIT_0A => X"A2020010100007865421432121804021C20452880C2D200000045C18C0E0000A",
INIT_0B => X"371097006026226495446E2110AE4417411204400000306B8186185C42900693",
INIT_0C => X"A00308003080030800308003080030800308001840018400400602A018809800",
INIT_0D => X"4008081010108003C000210020460801001FB3650C50DB13111C0D95C20C2030",
INIT_0E => X"14804032007E281F840C00284A17210001060D8306C18360C1380A0260CB9808",
INIT_0F => X"1555D5D79BBEF8E50B041029075982BF3873041029079982BF39748AA0AC8000",
INIT_10 => X"5156AEA479BFD7F7F3041029075982BF3E73041029079982BF3F632C5F96D3C1",
INIT_11 => X"932C5F96A595405FC7F1CFEBC7586C4100A53162B47FD7E39FFEECE159870234",
INIT_12 => X"39464006FE037ACFB88083A99E06271BB0CA207DFDD5920057E0B001B0EBCC79",
INIT_13 => X"6F5DF5CA2A002DD51B6F7FC4A411D1E8D44517F14EAFE36E55150016EA8DB73E",
INIT_14 => X"9DB84953C30351452A13D55CFFA76E928E3891F148B30399F5FB7F28C800DFA0",
INIT_15 => X"110155AC57DFEAEF1005475F1D1F608819CF0EE76E12C824ADD9089715F25FAF",
INIT_16 => X"0D8360D834041A41A0000010180C02801680460FC900052FA10DC0006DA4881C",
INIT_17 => X"D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D836",
INIT_18 => X"8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360",
INIT_19 => X"B000000000000000000000000020D8360D8360D8360D8360D8360D8360D8360D",
INIT_1A => X"1451451451448982C8A82E0820825942495377D9D701DC2E784601F8D187BEF8",
INIT_1B => X"4A2512A954AA5528944A25555145145145555555145145145555555145145145",
INIT_1C => X"FFC00000944A25128944A25128944A25128944A25128944A25128944A2512894",
INIT_1D => X"A5D2E820BA550000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFBFDFEFAAD142010007BEAB55FFAA821FFFFFFFFFFFFFFFFFFFFF7FBD74A",
INIT_1F => X"1FF002A821FFFFFFFFFEFF7D16AB55A2D542000A2D5400BA0800021FFFFFFFFF",
INIT_20 => X"DFFFFFFFC0010F7842AA10F780021FFFFFBFDF45A2D56AB45FFFFD54BAFF8000",
INIT_21 => X"6AB45A28000010082A975EFA2D140145007BC21FF5D2AAABFFF7D168B45AAD57",
INIT_22 => X"BC214555003DE10A2FBEAA00000002010552E95410AAFBD75FF5D7FEAB550051",
INIT_23 => X"04174AA5D00020BA555542145A284155FF5D517FE000004020AA552E80000F7F",
INIT_24 => X"00000000000017400082E954AA0800154AA0855575FFAAD57FE005D7BD740008",
INIT_25 => X"FFFFFDFEFF7FFD74AA552A820AA490A000000000000000000000000000000000",
INIT_26 => X"A080A051FFFFFFFFFEFF7F1FAFD7A2D5400001C7BEDB7DEBA4871FFFFFFFFFFF",
INIT_27 => X"6DFFFBD54AAE38E021FF0824821FFF7F1F8FC7EBD568B7DB6DF47000AADF400A",
INIT_28 => X"BC7E3D56AB7DB6DF78FD7EBF1C2000F78A2DA38E38A021C7E3F1F8F55AADB6FB",
INIT_29 => X"25EF497FEAB7D145B6FB45AA8E070281C20925FFBEDB451451C7BC01EF4124AD",
INIT_2A => X"00092412A87010E3F5C0145410E3DE28B6FFE8A101C0E05010412495428AAF1D",
INIT_2B => X"B7AE385D7FD74381400124825D0A000BA555F47145BE8A105EF555178E381C0A",
INIT_2C => X"00000000000000000000000000000154280024924AA1404174AA0055505EFBED",
INIT_2D => X"A80155FFFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA082A8000000000000000",
INIT_2E => X"F7FBD5410AAFBC00AA002A955FFF7FBFDFEFFFD568B45AAD5400005D7BFFFEFA",
INIT_2F => X"5AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF0000021EFF7D16AB55A2D56ABEF",
INIT_30 => X"45557BC21FF08003FF55AAD168BFFF7FFEAB45AAD140010F7AABFEBAAAAA8214",
INIT_31 => X"4100000154AAA2D1421FF007BE8BFF557BFDF55A2AA974AA5D04001EFFFFFD55",
INIT_32 => X"01EF55516AAAA5D2A82000082E95400A2D542155002ABDEBAF7FBE8A00552E95",
INIT_33 => X"174AA0855421FFFFFBEAAAA5D7BD74BA5D0002010552E820AA5D7BD7545F7AA8",
INIT_34 => X"0000000000000000000000000000000000000000000000174BA0004000AA5500",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000001000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000008128000000000000000000000024001620280000000000354200004008",
INIT_04 => X"000058800004C4024024001210001054B1C822009640000E2000002604003000",
INIT_05 => X"07008000E0200000000000000000200604000000001C04000026400000002C40",
INIT_06 => X"000000000000000004C010B35420015040000000002C42010010200004C83810",
INIT_07 => X"06E200201C00A14080082B26208008A009001201014022404402800408408020",
INIT_08 => X"00004180261C81210031000004340000200008105428020568040213003499C0",
INIT_09 => X"0000000990000000B0C308000000000860200160000000000038380000000000",
INIT_0A => X"10000000000005860000000080A0002060204080000000000004540800000000",
INIT_0B => X"00000000000000020001000022000000000000000000178000F8000101259000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000108000EC000000000000000010004B200000000000000000000000000",
INIT_0E => X"2000000000062801800400000000000000000000000000000000000000000000",
INIT_0F => X"828008084451B81A70AB3006BA0011400760AB3006BA0011400680F020968348",
INIT_10 => X"30B8011204082248A0AB3006BA0011400160AB3006BA0011400084C780687DBA",
INIT_11 => X"64C78068796E80A00802301BC0A7531EDD98E73B02800804620D030F873EB49F",
INIT_12 => X"B0A936B00000002044F091A860700FF9198AA115D5DA37F7A80C8A3604001C06",
INIT_13 => X"0000098551AC9000000000314E01F9F30198600631448410A2A8D64800000081",
INIT_14 => X"1046B2E00303842281C80A23004411AD661891F15148A4420804241526D60000",
INIT_15 => X"66A4A9D335F3D282000C6C5456C84850F61050C411AD6284FDA861682805A04A",
INIT_16 => X"0000000000000000000000000000000000004600C00138000030880042023043",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"9000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C30C30C30C3451046260A9A69A603924554117747E18E0218CC01400163A20C",
INIT_1B => X"26934984C26130984C26130C30C30C34D30C30C30C30C34D30C30C30C30C30C3",
INIT_1C => X"FFC000004C26130984C26130984C26130984C26130984C26130984C26130984C",
INIT_1D => X"A5D2A800105D2E80000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFF7FBD74AA5D2E820BA55003DFFFFFFFFFFFFFFFFFFFFFFFFFD54A",
INIT_1F => X"B55FFAABDFFFFFFFFFFFFFFFFFDFEFF7FFD54BA5D2EA8BFFFF84021FFFFFFFFF",
INIT_20 => X"8B55A2D540010007BEAABAA2AE821FFFFFFFFFFFFFFBFDFEFAAD142010007BEA",
INIT_21 => X"021FFFFFFFFFEFF7D16AB55A2D542000A2D5400BA08003DFFFFFFFFFFFFF7FBE",
INIT_22 => X"FD54BAFF80001FF002ABDFFFFFFFFDFEFA2D56AB45AAFBD74AAFFD5420100804",
INIT_23 => X"FBE8B45AAD568BFFF7FBD74BAFF802ABFFFFAE821FFFFFBFDF45A2D56AB45FFF",
INIT_24 => X"0000000000002ABFFF7D168B45AAD57DFFFFFFFC0010F7842AA10F780155FFF7",
INIT_25 => X"FFFFFFFFFFFFBD54AA5D2A80000412A800000000000000000000000000000000",
INIT_26 => X"7E384071FFFFFFFFFFFFFFFFDFEFF7FFD74AA552A820AA490A38FFFFFFFFFFFF",
INIT_27 => X"D7A2D5400001C7BEDB7DEBA4BAFFFFFFFFFFFFF7FBFDFD7EBF1D24AA5D2AADBD",
INIT_28 => X"FFFFFFBFDFC7E3F5EAB45AAD140000007FEFA92A2AA851FFFFFFFFFEFF7F1FAF",
INIT_29 => X"74AAE3DF400000004021FFF7F1F8FC7EBD568B7DB6DF47000AADF400AA080A3F",
INIT_2A => X"F8F55AADB6FB6DFFFBD54AAE38E021FF0824BDFEFE3F1F8FD7AAD16DB7DBEFBD",
INIT_2B => X"A2DA38E38A125C7E3F1EAB55B6DB6FBD7E3F5D04AAFF8A2DBD7E3A0821C7E3F1",
INIT_2C => X"000000000000000000000000000002DBC7E3D56AB7DB6DF78FD7EBF1C2000F78",
INIT_2D => X"82AA8BFFFFFFFFFFFFFFFFFFFFF7FBD54BA552A80010002A8000000000000000",
INIT_2E => X"A2D5400AA552ABDF55A280155FFFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA0",
INIT_2F => X"FF7FBFDFEFFFD568B45AAD5400005D7BFFFEFAA8028BFFFFFFFDFEFF7FFFFF55",
INIT_30 => X"10AAFBC00AA002ABDFEFF7FBFDF55AAD16AB55AAD140010007BFFE10AAAA955F",
INIT_31 => X"B45A2D57DFFFFFFFD54AAA2FBC20100800021EFF7D16AB55A2D56ABEFF7FBD54",
INIT_32 => X"FF45AA8002145AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF00003FFEFA2D56A",
INIT_33 => X"EAB45AAD140010F7AABFEBAAAAA82155AAD568B55FFFFFDF55A2D1400AAF7AAB",
INIT_34 => X"00000000000000000000000000000000000000000000003FF55AAD168BFFF7FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000002000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"000079800014CC02C034001600000000000000101EC0012EE0C0026E1E80F000",
INIT_05 => X"1F0FF433EFF0440C3902100002203F2EFC040388137C3E20C8EEC00284033CC0",
INIT_06 => X"7000660016490201700000000002FF57C8E8840155FDC0000010E40087D8787A",
INIT_07 => X"4000040007700000000000000001080FF900160000000200C00080001840BFE4",
INIT_08 => X"0009FFBFE5181606000410A4000004202AA8043E0000000000000001209244C0",
INIT_09 => X"0001227FB0000000F7DF78020004011FEFE00000000020031502000083880200",
INIT_0A => X"00000000000015BE0000004000000100000100506002008C2007D5FC80000024",
INIT_0B => X"0020000000000000000000000000000000210018800000000000000010000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000020",
INIT_0D => X"0008000000100000010000002000080101FFB600000000000000000000000000",
INIT_0E => X"0000003007FE29FF800C00000001002040000000000000020480002E42429C00",
INIT_0F => X"000000004D4E180010040000400000001E60040000400000001E6010003C0000",
INIT_10 => X"04000000000094B1E0040000400000001E60040000400000001E608040000004",
INIT_11 => X"0080400002000000000033628000100100000004000000006170C00080010000",
INIT_12 => X"B0020000000000295810000000A100020614148002000000000004307CC3CC00",
INIT_13 => X"000525802000000000014AC000120200000000003F0D800020100000000000A4",
INIT_14 => X"000020020C0C00000000002E2D000001006204040000000005786C0040000000",
INIT_15 => X"004000100A0C0939BEE1810080200000E0CE0EC000010020000000000000AE8A",
INIT_16 => X"000002008040400400C08080000000000049F6FFC01000000000000080080080",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"6902001000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"186186186190324C1090D0F3CF3CD039A060000600704000201120AB02090082",
INIT_1B => X"0C86432190C86432190C86596596596596596596596596596596596596596186",
INIT_1C => X"FFC00002190C86432190C86432190C86432190C86432190C86432190C8643219",
INIT_1D => X"A552A82010080400000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD54AA5D2A800105D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"0BA5500001FFFFFFFFFFFFFFFFFFFFFFFBD54BA552A8001000003DFFFFFFFFFF",
INIT_20 => X"FFEFF7FFD74BA552E801FF002E821FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E82",
INIT_21 => X"BDFFFFFFFFFFFFFFFFFDFEFF7FFD54BA5D2EA8BFFFF843FFFFFFFFFFFFFFFFFF",
INIT_22 => X"142010007BEAB55FFAA801FFFFFFFFFFFFFFBFDFEFFFD542000082EAAB55AAAA",
INIT_23 => X"FFFFFFFF7FBFDF55AAD140000087BE8B55F784021FFFFFFFFFFFFFFBFDFEFAAD",
INIT_24 => X"0000000000003DFFFFFFFFFFFFF7FBE8B55A2D540010007BEAABAA2AE975FFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA552A820001400000000000000000000000000000000000",
INIT_26 => X"81C0038FFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2A80000412ABFFFFFFFFFFFFF",
INIT_27 => X"EFF7FFD74AA552A820AA490A021FFFFFFFFFFFFFFFFFFEFF7FBD74BA5D2A8002",
INIT_28 => X"FFFFFFFFFFFFFFFBFDFEFFFFFD54BA5D2A801C7142E871FFFFFFFFFFFFFFFFDF",
INIT_29 => X"0010142AAFB7DBEAEBAFFFFFFFFFFFFF7FBFDFD7EBF1D24AA5D2AADBD7E38438",
INIT_2A => X"FFFEFF7F1FAFD7A2D5400001C7BEDB7DEBA4871FFFFFFFFFEFF7FBF8FD7E3D14",
INIT_2B => X"FEFA92A2AA925FFFFFFFDFEFE3F1FAF45A2D142010087FEDB55F78A051FFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFBFDFC7E3F5EAB45AAD140000007",
INIT_2D => X"02ABFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005D040000000000000000",
INIT_2E => X"F7FFD74AA5D2A800BA550428BFFFFFFFFFFFFFFFFFFFFF7FBD54BA552A800100",
INIT_2F => X"FFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA082A821FFFFFFFFFFFFFFBFDFEF",
INIT_30 => X"AA552ABDF55A2802ABFFFFFFFFFEFF7FBFFFFFF7FBD74BA552A80145552E955F",
INIT_31 => X"FEFF7FFEAB45AAD1420105D2ABFFFFFFAEA8BFFFFFFFDFEFF7FFFFF55A2D5400",
INIT_32 => X"DF55F7AE955FFF7FBFDFEFFFD568B45AAD5400005D7BFFFEFAA80175FFFFFBFD",
INIT_33 => X"6AB55AAD140010007BFFE10AAAA821EFF7FBFDFFFAAD168B55A2D542010007BF",
INIT_34 => X"00000000000000000000000000000000000000000000003DFEFF7FBFDF55AAD1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"084A76341244919000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"000079800014CC03C075161E001118653D2408041FC004AEF000816E1C11F541",
INIT_05 => X"3F0F807BFFE000240100004683103E7FFE02482553FC3C0204EFC25010143CC0",
INIT_06 => X"1100441004201014B1709C910102FF5FC0A0000101FFE4036450E08247F87870",
INIT_07 => X"08750504800680102542AD800504530FF9061E8026998E9A00402CC25BD0FFFC",
INIT_08 => X"0011FBFFE04691A5A00101818A6800088228000001A044C8168480D010F200AA",
INIT_09 => X"B6E85A7FF080AC70FFDF78220010841EFFE7116E144071268DFD3E4C24040100",
INIT_0A => X"3151518A8A31B7FE00040009814C089202225412115428C03BC7D7FC15025B1A",
INIT_0B => X"1B1883007104032901CC63410ABD249C4B338934404037FC8BFE18008083B444",
INIT_0C => X"D9228D9228D9228D9228D9228D9228D9228D99146C9146C84006309044081A00",
INIT_0D => X"48000201800500941044312000900D4621FFBE00080081529904595123203040",
INIT_0E => X"308162029FFEADFF8050250010030165290008800440022201082401A002000C",
INIT_0F => X"5001318048A004A6C0D2820302C005A83480D1820302A009B02B101390C0CB28",
INIT_10 => X"485101408904831400D1820302C005A83480D2820302A009B02B021A85C09411",
INIT_11 => X"FA1A85C08834600024D052C1051E0B92D400360520202682C19024B6164E3004",
INIT_12 => X"C1B0D6404093E22A2012418A9D1D44ADD9E0F174103820101C0B8160D5516259",
INIT_13 => X"6C88660D8AA288209E615100280DA0052000C5006402000206C55144104D510C",
INIT_14 => X"024500A0D50020C04023033C52009144231D902818100C90058010361AC80812",
INIT_15 => X"198A12202386454988140600C0181500A13E830011008B0374007000B4E0CD00",
INIT_16 => X"008020080224004002000000703804008001F7FFF01B982B01258088C008CC41",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"F000000000000000000000000020080200802008020080200802008020080200",
INIT_1A => X"7DF7DF7DF7DFFFFEFEFFFE79E79FFFF3BC1FF3FDDFEFFFBEFFE7DF84081EFEFB",
INIT_1B => X"FEFF7FBFDFEFF7FBFDFEFF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF",
INIT_1C => X"FFC00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"A5D2E80010000400000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA552A8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"0105D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E80010552EBFFFFFFFFFFF",
INIT_20 => X"FFFFFFFBD54BA5D2E82010002ABDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A80",
INIT_21 => X"001FFFFFFFFFFFFFFFFFFFFFFFBD54BA552A800100000001FFFFFFFFFFFFFFFF",
INIT_22 => X"BD74AA5D2E820BA5500001FFFFFFFFFFFFFFFFFFFFF7FBD74BA5D2E800BA5D00",
INIT_23 => X"FFFFFFFFFFFFFFEFF7FBD74AA552A800BA5D2E821FFFFFFFFFFFFFFFFFFFFF7F",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFEFF7FFD74BA552E801FF002E975FFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E800000800000000000000000000000000000000000",
INIT_26 => X"05D2ABFFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8200014003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFBD54AA5D2A80000412ABDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2E8000",
INIT_28 => X"1FFFFFFFFFFFFFFFFFFFFF7FBD54BA552E82028002AB8FFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74AA5D2E800AA5500021FFFFFFFFFFFFFFFFFFEFF7FBD74BA5D2A800281C0000",
INIT_2A => X"FFFFFFFFFFDFEFF7FFD74AA552A820AA490A071FFFFFFFFFFFFFFFFFFEFF7FBD",
INIT_2B => X"A801C7142E955FFFFFFFFFFFFFFFFDFEFF7FFD54BA5D2E80082492E871FFFFFF",
INIT_2C => X"0000000000000000000000000000038FFFFFFFFFFFFFFFBFDFEFFFFFD54BA5D2",
INIT_2D => X"D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008000000000000000000",
INIT_2E => X"FFFBD54AA5D2E800005D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF7FBD54BA552A80010002ABDFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"AA5D2A800BA5504021FFFFFFFFFFFFFFFFDFEFF7FBD74AA552E820BA002AA8BF",
INIT_31 => X"FFFFFFBFDFEFFFFFD54BA552E800BA5D04021FFFFFFFFFFFFFFBFDFEFF7FFD74",
INIT_32 => X"0000082A955FFFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA082A955FFFFFFFF",
INIT_33 => X"FFFFFF7FBD74BA552A80145552E975FFFFFFFFFEFF7FBFDFFFFFFBD74AA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000002ABFFFFFFFFFEFF7FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"431965109E4481D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"492C0020220001010E4916C884DCD607E5EC2A344103E48003D0800023D0072C",
INIT_05 => X"00107C441001100D620A06D683018001023D37E5088043620101179092540112",
INIT_06 => X"401002010042384D223C19C3552800081ADA0E054402365774611E047020008E",
INIT_07 => X"491EC04ED017AB5497EB923F08182E20020689B735011FBFE7BC062602944019",
INIT_08 => X"154A00401D4425ADA9035BE19C8F9442A8801200F4C9D7AC8093A051727B2AC3",
INIT_09 => X"9A50020040E48D50080002B00A0C00801014541E9504703680017F6CB4050700",
INIT_0A => X"8151538A8A738041C23020131A80CFDFF3FE509A907C6AC05040220409009031",
INIT_0B => X"2D040050110081E9528963546278008AA80381B4000500026800000109379864",
INIT_0C => X"1C2A81C2A81C2A81C2A81C2A81C2A81C2A81C9540E1540E00140000610000320",
INIT_0D => X"594A06870A9CA0D458D131652A154D46B6000850800801628013456520CA0928",
INIT_0E => X"02080448C00044000A1EC1C44140D101A54280A14050A028500A84F02842A24C",
INIT_0F => X"0061338359E0C4E6C256690581800F1C3E82562B0581200F1C3F081456022804",
INIT_10 => X"2C438100AB8581B602562B0581800F1C3E8256690581200F1C3F1238473F1210",
INIT_11 => X"2238473F0E1050083750B3E4275F829547008600C030374361FA2CEE046D4812",
INIT_12 => X"C1128C4CC012A66F61154C019511628756231018500C00203E13806156516078",
INIT_13 => X"54CDE608AA612C0096C37B00D1724801A0009C606D1221D104553096004B61BC",
INIT_14 => X"870B012A41E0F0600035842E7601C2C4AC68A98810080AA825A8902251899802",
INIT_15 => X"58234A89637E00D0A1080301401C390320188321C2C0B13890105800D520AF94",
INIT_16 => X"8822088222F110111B281A54753AA004002601001918008C10912A4440B24E8B",
INIT_17 => X"8220882208822088220882208822088220882208822088220882208822088220",
INIT_18 => X"2008020080200802008020080200802008020080200802008022088220882208",
INIT_19 => X"E82891448000000001FFFFFFFFC8020080200802008020080200802008020080",
INIT_1A => X"3CF3CF3CF3DFFBFEFEBEEEFBEFBEFBEBFDF7F7FBDFD1FE3EFBD7ADFBF7EFBEFB",
INIT_1B => X"FE7F3F9FCFE7F3F9FCFE7F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"FFC00001FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"A5D2E82000000000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8000008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74AA552E8000055003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A82",
INIT_21 => X"BFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E80010552EBFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD54AA5D2A800105D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A82000552A",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD54AA5D2A800005D2EBDFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000000001FFFFFFFFFFFFFFFFFFFFFFFBD54BA5D2E82010002AA8BFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100004000000000000000000000000000000000",
INIT_26 => X"008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA552A8200014003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E800105D043FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"54AA5D2A82010552EBDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2E800005D2ABF",
INIT_2A => X"FFFFFFFFFFFFFFFFFBD54AA5D2A80000412AB8FFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E82028002AA8BFFFFFFFFFFFFFFFFFFFFFFFBD54BA552E80038492EB8FFFFFFF",
INIT_2C => X"00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFF7FBD54BA552",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000040000000000000000",
INIT_2E => X"FFFFD74BA552A8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E800000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005D043FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"AA5D2E800005D2EBDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA552E8001055003FFF",
INIT_31 => X"FFFFFFFFFFFFF7FBD54BA5D2A820105D2ABDFFFFFFFFFFFFFFFFFFFFFFFFBD54",
INIT_32 => X"00AA082EA8BFFFFFFFFFFFFFFFFFFFFF7FBD54BA552A80010002AA8BFFFFFFFF",
INIT_33 => X"FDFEFF7FBD74AA552E820BA002AAABFFFFFFFFFFFFFFFFFFEFF7FBD74BA552E8",
INIT_34 => X"0000000000000000000000000000000000000000000000021FFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"2C4360101A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"00017B810015DC03D034201E14000036486008101FC0002EE006297E1C05F561",
INIT_05 => X"BF0F817FFFE80100004044800080BEFFFC0248005FFC3C18A5FFC2444484BCC0",
INIT_06 => X"B0801408110000109127E0500002FFDFC000000001FFC0832050E00047F97870",
INIT_07 => X"00D1D72040048D00388387D03D0E591FFD201F862691DFBE077C2BC45B40FFE4",
INIT_08 => X"001FFBFFEC440501A5604B31062356282AA84200D12342113EDC400000045828",
INIT_09 => X"25A890FFF0002023FFDF79000000000EFFE309606020008005FC000000402000",
INIT_0A => X"30000000000037FF50010103134CAFDF03BA18000F39A0106F87D7FA84024B02",
INIT_0B => X"1B188300624483890564084198AD249C43300C00415037FC83FE1840C0902400",
INIT_0C => X"C1010C1010C1010C1010C1010C1010C1010C10086080860840063090442A1800",
INIT_0D => X"0001403000100200180480000095280001FFBF040C40C81119A41C1443243050",
INIT_0E => X"32A163821FFEAFFF805025E00853B92588000400020001000020A80180080020",
INIT_0F => X"90401486148484054395E27E428002A4200397E07E422002A420100382FCC308",
INIT_10 => X"641100C0788417000397E07E428002A4200395E27E422002A420110A51C01C05",
INIT_11 => X"C90A51C01A2490040590C08120558C1759BE1C05A0400383808800DA1929F728",
INIT_12 => X"00CE720000136006000215EA0A4833A32C8832050028603050014031B3950000",
INIT_13 => X"6C00C006658280009A2030108B14AC05C00112405222088B8332C140004D1018",
INIT_14 => X"A2659196B6808060201281004228996085F10020180C030880D11019CE400002",
INIT_15 => X"0108152A49DC7143F01C04240030720641E0A028996483A17204680410A04104",
INIT_16 => X"040100401000080080000000000002001201F7FFC0011C2F81A48080CA32800A",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_19 => X"0000000000000000000000000000401004010040100401004010040100401004",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000020000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFC0000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2A8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E80",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8000008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA552A8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A820000004",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA552A8201000043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E8000055003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA552A8200008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001008043F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA552A8200014003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E800105D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E820101C003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552",
INIT_2D => X"0043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA552A8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001008043FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74AA552A8200008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"200055043FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005D043FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD54AA552E8001055003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA552E8",
INIT_34 => X"00000000000000000000000000000000000000000000003DFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"00003A2E200811000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"000079800014CC03C034001E04010850300000101FC0002EE000006E1C00F500",
INIT_05 => X"1F0F8033FFE000000000000000003E2FFC024800137C3C0000EFC00000003CC0",
INIT_06 => X"000000000000000091C115500002FF5FC000000001FFC0000010E00007F87870",
INIT_07 => X"10E600084002040A10812A000500590FF9001F95406A8000037230C01840FFE0",
INIT_08 => X"0001FBFFEC4695A501604A000C7585080002C200408102F16C0184800026C92C",
INIT_09 => X"24A8107FF0000000FFDF78000000000EFFE001600000000005FC000000000000",
INIT_0A => X"30000000000037FF4000000AA0354000019C4000012800002387D7F804024B02",
INIT_0B => X"1218830060040A04000400000801241443300800404037E883FE180000000000",
INIT_0C => X"C1000C1000C1000C1000C1000C1000C1000C1000608006084006301044081800",
INIT_0D => X"00000004800B0000000000000000000001FFBE00080080101904181003003000",
INIT_0E => X"B08062021FFEADFF800020800000002088000000000000000000200180000000",
INIT_0F => X"D0210840009181008024A00043601100210024A00043C0110020901382CCCB28",
INIT_10 => X"0C920180040A03080024A00043601100210024A00043C01100209240C840C201",
INIT_11 => X"1A40C840A604E0080820009908008341B000A821207008200289001006832086",
INIT_12 => X"0166B40600800082041205EC00044C1ACB66C37542082030281E058000101281",
INIT_13 => X"0010480B27A004300004103160DB3005E000618040C022000593D00218000209",
INIT_14 => X"880012BBFF20406040084210C062000C2A2DDD00180C04504086002CD680C010",
INIT_15 => X"4106020804295C98F80400008040CC0582169022000C2876C404780028500160",
INIT_16 => X"000000000000000000000000000000000001F7FFC001B823018F008800088052",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"C800000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"7CF7CF7CF7D933CC3090CABAEBAFF969319815DD5EDCF9822659AE7B095A220C",
INIT_1B => X"1E0F0783C1E0F0783C1E0F7DF7DF7DF3CF3CF3CF3CF3CF7DF7DF7DF7DF7DF7CF",
INIT_1C => X"FFC000003C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C",
INIT_1D => X"A5D2E82010080400000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"00000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E800000800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8001000003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100804000000000000000000000000000000000",
INIT_26 => X"000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"A8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000043FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008040000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8000008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"000008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2A8001008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00002000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"924279824C94CC1BE0B4001F20000000020380401FE0082EF000106E1C00F500",
INIT_05 => X"1F0F8033FFF048202582800100523E2FFE024820137C3C0040EFE02000003CE4",
INIT_06 => X"F10466105670019C900000100002FF5FC0E0801101FFC0000010E08A07FC7870",
INIT_07 => X"0000040000000000000000000500590FF9001F0000000000033020C01840FFFC",
INIT_08 => X"0001FBFFFD0004000100502000011400000282004001020000000001009015C0",
INIT_09 => X"2CB8DA7FF8004000FFDF7C062031863EFFF75D78004001010DFC000020050100",
INIT_0A => X"30000000000037FFC00602000000000001980400002800032387D7FE94FBEF2B",
INIT_0B => X"9258830060040200000400000801243443B00808404037E883FE180C00000000",
INIT_0C => X"C1000C1000C1000C1000C1000C1000C1000C10006080060840077330C4889CC2",
INIT_0D => X"0000000000000000000000000001280001FFBE00080080101904189003003000",
INIT_0E => X"30A063021FFEADFF805025C0304001E58906088304418222C108A009A0904000",
INIT_0F => X"1000000000100100000480000200100000000480000200100000100380F0C308",
INIT_10 => X"0010000000080000000480000200100000000480000200100000000040400000",
INIT_11 => X"0000404000040000000000080800000110000000200000000200000000012000",
INIT_12 => X"00021000000000800002018C0100000208000008001220000000040040000080",
INIT_13 => X"0010000020800000000400000010200200000000008002000010400000000200",
INIT_14 => X"0800000210000080010000008002000000210000201000000002000042000000",
INIT_15 => X"0184000000084000000006050000000002000002000000204000000000000020",
INIT_16 => X"08822288226410410346010000000400A011F7FFE00318230104008000008000",
INIT_17 => X"8822088220882208822088220882208822088220882208822088220882208822",
INIT_18 => X"8220882208822088220882208822088220882208822088220882208822088220",
INIT_19 => X"0404000017FFFFFFFFFFFFFFFFE0882208822088220882208822088220882208",
INIT_1A => X"492082492085048029890AD34D35FDD04A165129432D518B45265EFC30760AED",
INIT_1B => X"C46231188C46231188C462492492492492492492492492082082082082082082",
INIT_1C => X"FFC000058AC562B158AC562B158AC562B158AC562B158AC562B158AC562B158A",
INIT_1D => X"A5D2E820100800000000000000000000000000000000000000000000000003FF",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100000",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000043FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"4A53D958C50000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"DBFAFBD7FB1CDEBEF1BE17F7AC88042787FBFFF8FEE9FF7EE6F4C0EE1FFAF869",
INIT_05 => X"5F0FFEB3EFFEFFBDA7F7FED508707E2EFEBF6FFEB37C3FF302EEEDFF9B487CF6",
INIT_06 => X"74EADE4EBDFDAC9930F6F8129E3FFFF7C3E3A74667FDDB7FB870FF30FFDEF87F",
INIT_07 => X"8173840C07783060C72DF7D828912E6FFB80162776F3BFB7077E82255E40BFEF",
INIT_08 => X"4769FFBFE43C872321367036163F1C0820A3063F460D1AEFC000060042648C41",
INIT_09 => X"BEFB967FBD13D981F7DF7D7E6171AF3FEFE8A3E679FAC1FD1FFFBEB000763A84",
INIT_0A => X"F3A3AD1D1DAD7FBE7D67D7F3BB79CFFB83BF14EC1E7D7300B017F5FFE6FBEF73",
INIT_0B => X"52199F58F6EE6F5E7FAC4C03DB856CD4CF720FE8C4427FF8CFFE38FF7F6BD928",
INIT_0C => X"F78C0D78C0D78C0D78C0D78C0D78C0D78C0D7A606BC606B8C56F7730ECCDBDF1",
INIT_0D => X"EA035CF6100C0E60FB9FC3A80EF69A04DFFFF7FF5E75FF341B867D3683A03A40",
INIT_0E => X"36B867027FFFF9FF8FAFAA3ADEBFB9726BAF5FD7AFEBD7F7EFFD7ACDB7F947F0",
INIT_0F => X"10003E020080A40403E8BD8002000FC02003E8BD8002000FC02010979AFFE36C",
INIT_10 => X"80100000EE00034003E8BD8002000FC02003E8BD8002000FC020037B0040A000",
INIT_11 => X"037B0040C00400003D80008160400FD81341C00020003B80008C00801EF02853",
INIT_12 => X"01F1190981038406809677FA080468C46A81080581002000780C8001C8100201",
INIT_13 => X"7080D00F90D162001C803411FC0024080001F80040026C0807C868B1000E401A",
INIT_14 => X"B02013F810503A00003E020042AC080CEB01228A80000F600080123E23213040",
INIT_15 => X"61F810087520750001064180807868000110C02C080CFA0042400000F8800105",
INIT_16 => X"5FD7F7FDFF7EFEEFF3EEC3FF7FBFFBCB7FFFFEFFE00BFF7FEBF420800EC0CBEE",
INIT_17 => X"FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F",
INIT_18 => X"D7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5",
INIT_19 => X"6DAE443237FFFFFFFFFFFFFFFFF5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5F",
INIT_1A => X"4D34D30C30DD795EAA6AFC38E38EA3AB788962B79E923C2CD990A7D3B4A9FC37",
INIT_1B => X"26130984C26130984C26130C30C30C30C30C30C30C30C30C30C30C30C30C30C3",
INIT_1C => X"FFC000004C26130984C26130984C26130984C26130984C26130984C26130984C",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"0842D85841000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"DBEAE5D6D91C2EBCE1B21EA72C00000007FBE7C8F8E9EF79E6D440E91FDAE061",
INIT_05 => X"5C8FFCB38FF6B68984B5BCE408347E28FEBF6FEEB3723F7102E8EDBF8A4872F6",
INIT_06 => X"946ACF46ACE0841A00006A089E3FFF27C3032646EFF1DB7FA868FE30EF1CE47E",
INIT_07 => X"8000000A20083060C00C81882A008C6FF880060424B39FB6037F00051C003FE0",
INIT_08 => X"4761FA3FE4010440410844060001040A00002200460D1A060000050400000010",
INIT_09 => X"FEEB027E390A4881C7BEFC5F6171CE2F8FE823E778DAC16C1FFBBC9000315895",
INIT_0A => X"F606013030213C3E2D62D6E21259CFDB039E806C024531008017C1F826FFEF41",
INIT_0B => X"5219AB5AF86F7D5E382A440349816DD4C7560B60D4427FF0C7FEBABF3F6BD108",
INIT_0C => X"E3440C3440C3440C3440C3440C3440C3440C3C2061A2061AD46FF730E5CCBCD5",
INIT_0D => X"6203E8FC10080A20ED1D41880CC61A044DFFC6EB5AB5B7941BC63F1683803C00",
INIT_0E => X"B88572023FFE91FF98AEAA1AC6AC9A3A4AAD5B56ADAB56D5AFD572C597B14750",
INIT_0F => X"10003E020000260403C8948002000EC0000BC8948002000EC00010878AC3CB8A",
INIT_10 => X"80100000EE0000400BC8948002000EC0000BC8948002000EC000097B00402000",
INIT_11 => X"017B0040400400003D80000070400DD81041400020003B80000410801AF02041",
INIT_12 => X"05D11101010384008086378A080428C46A80080081002000780C800188000301",
INIT_13 => X"7080102E909042001C800409FC0020080001F80000007C0807484821000E4002",
INIT_14 => X"F02003F810100A00003E020000BC0808EB01020280000F60000002BA22202040",
INIT_15 => X"21F810007520750000024080807868000100403C0808FA0040400000F8800001",
INIT_16 => X"5B56D5B5EF3AF6AF6389C2FE128971AB2DDDF8FFE0031B776BF4208006C0C926",
INIT_17 => X"B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D",
INIT_18 => X"56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5",
INIT_19 => X"238B443A3FFFFFFFFFFFFFFFFFD5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B",
INIT_1A => X"00000000000F0080397908000000A4805F09C42D0200903950C086D420010825",
INIT_1B => X"8040201008040201008040000000000000000000000000000000000000000410",
INIT_1C => X"FFC00005028140A05028140A05028140A05028140A05028140A05028140A0502",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100804",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"461080404900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"00800040110102000902002000888400081045A8A00003C00000500000080008",
INIT_05 => X"0000000000024CA0A0101800032000400000000B800000014000000B08180000",
INIT_06 => X"0020280202802C00020800008A14002011110012220009A88800009A88000000",
INIT_07 => X"8108044200091224484510201000204000800020410000000080000104000009",
INIT_08 => X"132800000140200808021006108010422AAA8000224489028492201140092240",
INIT_09 => X"0001C800004080A0000002480B04008100011000088800081002C19020150B00",
INIT_0A => X"4353529A9A528000040040702080000000400064080011001050000200000018",
INIT_0B => X"01400048012220122A0004168110400004000040811600000400001036584108",
INIT_0C => X"36050160501605016050160501605016050160280B0280B00120008430660210",
INIT_0D => X"2A000C4210040860B188C0A8065302005A0040390010120500002002C0040010",
INIT_0E => X"8221050060001000028000080205001066000100008000400490020402010530",
INIT_0F => X"000000000000A00000081480000001400000081480000001400000800C010820",
INIT_10 => X"8000000000000240000814800000014000000814800000014000000100002000",
INIT_11 => X"000100004000000000000001400000080041400000000000000C000000100041",
INIT_12 => X"000101010100000480802A400000004000000800810000000000000048000000",
INIT_13 => X"0000900010104200000024000400000800000000000244000008082100000012",
INIT_14 => X"1000004000100A00000000000284000040000202800000000000120020202040",
INIT_15 => X"2050000010000000000240800000000000104004000040000040000000000005",
INIT_16 => X"010040108408420430E699AA42A1508104EA08000000810020000000044001AC",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"0506117080000000000000000000100401004010040100401004010040100401",
INIT_1A => X"4104104104006C1A8283AC618618EF10C0422205822140048D2E581E80DEC4D2",
INIT_1B => X"C06030180C06030180C060410410410410410410410410410410410410410410",
INIT_1C => X"FFC0000582C160B0582C160B0582C160B0582C160B0582C160B0582C160B0582",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0401D940CD0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"49B87A417315D20A313E17F1800000058013DDF8BE21F36E02F0D06E03E8F800",
INIT_05 => X"1F007E33E01A4D9C87525E5101603E6E023D27DA937C03E340EE25CB9B483C12",
INIT_06 => X"F0A05A0A15AD0C0130F6F0128A16FFF001E1870223FC3BFC98101F109FC6780F",
INIT_07 => X"8073800407781020476467D008910A4FFB80100332D1AE93059282215E408006",
INIT_08 => X"0221FF80003C832320342036063F08000001063F42050AEB4000221000248C01",
INIT_09 => X"9A51547F8C1111A0F041056A0100A11FE000916249A800B915FE82B020522900",
INIT_0A => X"42A2AD1515AD5780540541619968C76980E914E4163D53002017F405C409A42A",
INIT_0B => X"0140140816A22B126DA40C03531440800C2005C8800217F80C000055FF7C4928",
INIT_0C => X"268D0068D0068D0068D0068D0068D0068D006A68034680300021410028450530",
INIT_0D => X"AA01587410080C60AB0F42A804628200DBFFF13D04505B2500806522C0A40A50",
INIT_0E => X"941922006FFFF8000F8F80281A16A1504302058102C0816244B82A0CA25907D0",
INIT_0F => X"000000000080A40000283D80000001402000283D80000001402010901A7D6944",
INIT_10 => X"800000000000034000283D80000001402000283D80000001402002010000A000",
INIT_11 => X"02010000C000000000000081600002080341C00000000000008C000004100853",
INIT_12 => X"0021090981000006809076B20000404000010805810000000000000048100200",
INIT_13 => X"0000D0011051620000003410040004080000000040026C00008828B10000001A",
INIT_14 => X"B000104000503A000000000042AC00044000228A800000000080120421213040",
INIT_15 => X"607800081000000001064180000000000010C02C000440000240000000000105",
INIT_16 => X"05816258964C4A44A0C689FF3F9FFEC5D6DBFE0020096528A0B000000CC043EC",
INIT_17 => X"5816058160581605816058160581605816058160581605816058160581605816",
INIT_18 => X"8160581605816058160581605816058160581605816058160581605816058160",
INIT_19 => X"F506003017FFFFFFFFFFFFFFFFE0581605816058160581605816058160581605",
INIT_1A => X"5D75D75D75DFFFFEFCFDF7FFFFFF5DE7FC3DF3F2DDCFFFBEFFCF1F84421FFEFF",
INIT_1B => X"EFF7FBFDFEFF7FBFDFEFF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF75D7",
INIT_1C => X"FFC00007DFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDF",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"E800000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"3CF3CF3CF3DD7FDEBAFAFEFBEFBFFBFBB9DFF7FFDFF3FC3EFFF7FDFBBDFFFEFF",
INIT_1B => X"FE7F3F9FCFE7F3F9FCFE7F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"FFC00001FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"08425818000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"DB6A618248140C18E0B016872400000007EBA24058E1ECA8E2D400681FD0E061",
INIT_05 => X"1C0FFC338FF01009048084C400103E28FE3F6FE513703F7000E8E5B4825030F6",
INIT_06 => X"100046000460001800006800142AFF07C202060445F1F2572060FE82671C607E",
INIT_07 => X"00000008800020408008818838000C2FF800060424B39FB6037E000418003FE0",
INIT_08 => X"0441FA3FE4000400010040000001040880000200440912040000040000000000",
INIT_09 => X"BEE8027E38004801C79E7C162231862E8FE00166704041240DF93D0000000000",
INIT_0A => X"B00000000000343E002202021259CFDB039E0008024520000047C1F804FBEF01",
INIT_0B => X"121883107044094C1028400548812494C3120920404437F0C3FE180D89279000",
INIT_0C => X"C1000C1000C1000C1000C1000C1000C1000C18006080060840477330C4889CC0",
INIT_0D => X"400340B400080200481501000884080405FF86400800811019861D1403803800",
INIT_0E => X"308062021FFE81FF880EA000400098200C04080204010200810020C180904240",
INIT_0F => X"10003E020000040403C0800002000E800003C0800002000E8000100780C2C308",
INIT_10 => X"00100000EE00000003C0800002000E800003C0800002000E8000017A00400000",
INIT_11 => X"017A0040000400003D80000020400DD01000000020003B80000000801AE02000",
INIT_12 => X"01D01000000384000006118A080428846A80000000002000780C800180000201",
INIT_13 => X"7080000E808000001C800001F80020000001F8000000280807404000000E4000",
INIT_14 => X"A02003B810000000003E020000280808AB01000000000F600000003A02000000",
INIT_15 => X"01A81000652075000000000080786800010000280808BA0040000000F8800000",
INIT_16 => X"08020080223010010308025410082404A015F0FFE003182701B420800280C802",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_18 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_19 => X"0008004017FFFFFFFFFFFFFFFFC0802008020080200802008020080200802008",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFC0000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749803",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"441406267B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"0005802424830120024121209088809DF81454ACA01E03501D0A3B91E00F0A00",
INIT_05 => X"E0F001CC00012034C20B0232838F80D001C0100AEC83C008EF101A034C8CC300",
INIT_06 => X"2F1620F1721BA346AA2C95C5CB1400000161F84322000DA8C40F003C80030780",
INIT_07 => X"5939F36677EE1C387777622717EF711004A6818111086008E080FDC305940018",
INIT_08 => X"13160400195E83A3A0F61BC3929ECB622AABF5FF83860CEB164833F179B48CEE",
INIT_09 => X"01036D8004FDB47600000229410C61010016DC998C84B0128202C0DCB48F05D5",
INIT_0A => X"4400402A0A37000182502440888420247041E876810099D35F900002DB00105C",
INIT_0B => X"AD4434020CA2E0B32B01A752B078412A24818094151348062400E2A034D86444",
INIT_0C => X"3E2781EA781E2781EA781E2781EA781E2781C33C0613C0E21028840239452116",
INIT_0D => X"394818429A95E954868AD0E52273F54258000080808900C3807122C3E04E0338",
INIT_0E => X"8E3B15C94001120055704DC4A1624487E2489024481224091282C4300942A194",
INIT_0F => X"C06101C55D65C3E3F01F52FFC1E0013C1F801F52FFC1E0013C1F8090423D38A1",
INIT_10 => X"ECC381C0118796BE001F567FC1E0013C1F801F567FC1E0013C1F9085DFBF7E15",
INIT_11 => X"F885DFBF7E30F00C0270F3751F1FD00FECBF7E25C0700463E17B2C7F811FD7AD",
INIT_12 => X"C40FE6474190626D6491063597F9177B956EF378D33E4030061341F077C571F8",
INIT_13 => X"0C4DAE207F328E3082636B2807FFD80FE00007E03F7207D3E03F9167184131B5",
INIT_14 => X"1F4FE047EFA0CAE06101C53E3647D3F144FCDD22B81C0098E57D9081FCE8C852",
INIT_15 => X"38574FF31ADF08DBF81846A540049707E0FE3307D3F141FFB45478040570EED4",
INIT_16 => X"90240902C189601208A1102B4AA5584B4068000019A80098120BCA4C617635C9",
INIT_17 => X"0240902409024090240902409024090240902409024090240902409024090240",
INIT_18 => X"2409024090240902409024090240902409024090240902409024090240902409",
INIT_19 => X"9AA09426A8000000000000000009024090240902409024090240902409024090",
INIT_1A => X"104104104104431042720EE38E38AAF9A93E7131C136AD8E9B562CF03B2E8E78",
INIT_1B => X"F87C3E1F0F87C3E1F0F87C104104104104104104104104104104104104104104",
INIT_1C => X"FFC00001F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0",
INIT_1D => X"AAAAABDEBAF7AE8000000000000000000000000000000000000000000000C200",
INIT_1E => X"EFF7D142145A2AE800BA08514214555517DEAA5D7BFFEAAF7803FEBAF7FFD74B",
INIT_1F => X"E00A2FBD75FFFF84001550851555FF55517FE000055421FF00557DF45A2D5401",
INIT_20 => X"74BA552EBDFFF0004020005D5555555A2AABFFFF5D516AA00A28028A00AAAEBF",
INIT_21 => X"3FEBA082ABFE10AAAEA8ABA55517FF45A2AEBDEBAAAAAA8BFFF7D140010FF841",
INIT_22 => X"FD75FF0051401FF5D00154105504000BA5D2E97545A28028B450855401450804",
INIT_23 => X"FBFFF45A2FFFDE00002E801FFA2AABFE00FFFFD74AA085540000002E801FF557",
INIT_24 => X"0000000000002ABEFAA80001EFF7FFC20BAF7D1575450800020BA08517FF45F7",
INIT_25 => X"57803AEBAF7F5D74AAA2A03AA38BF8FC00000000000000000000000000000000",
INIT_26 => X"7A3F00516DA2D5451D7EBDB47155BC2A87092AAFA9257F1C5BC00AA5D7FF8EAA",
INIT_27 => X"00EA8000150A801C01C7142EBFBC7EB8005B55A85B555EF095F50578085BE8FC",
INIT_28 => X"BEAE3D542A004380124921D20975FFAAA1521FF492BF8F40B6AAB84AF555168A",
INIT_29 => X"8F6DE05B40480557A95A3A1C2EBAE28168ABAA2D43D568BC5400168E90E2F412",
INIT_2A => X"47B50A80095178157FEFA0742FA3AA28EA8168A954100071D2E90A855C7A00A3",
INIT_2B => X"0A8F57F6DA971F8F7FFFA42D16D1EAE925EA0BFEBF4AA09217F4905684170851",
INIT_2C => X"000000000000000000000000000002D57AAA8402A8743DBD202DA95568A95E80",
INIT_2D => X"17D34ABA5D7BEAAAAD786BCEAAFFD1564BA2282BFA02A2C28000000000000000",
INIT_2E => X"007F8B2B2D97D483AFA7BD9F5EFA87F57555AAFBD7555FFAE95408A8FDC31AD0",
INIT_2F => X"0A6AEA8FAF0451CA001D4845C2087383F79A5046A37B55F38415555797D63BFF",
INIT_30 => X"A7D7463CC508D07577BAFBD542000D382964A92B401E71D7581C33172EC0A030",
INIT_31 => X"0502828811FCD4EABDB1DFDFC8365A2FD5E04AA5780A8AAAD7AC3CA02003BEBB",
INIT_32 => X"4FF72AAADF245595157050790621F562B1122DA70C3808458881056A5502AA15",
INIT_33 => X"F6A03D4BFB79AFA4C5CB5F5896D55BBAAC55EAFAF86D35E4A92B4460D1506037",
INIT_34 => X"FC0000007FC0000007FC0000007FC0000007FC0000007FC07AAF12E00505D3FD",
INIT_35 => X"7FC0000007FC0000007FC0000007FC0000007FC0000007FC0000007FC0000007",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000400000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"650C00000848A0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000004208B00200E010800006667BE7000102C00080000040012010000080C",
INIT_05 => X"0080000000002020600100208D04414000800000000200004800080000800200",
INIT_06 => X"04022140220932C2038900000100000008082010000000800488000000020400",
INIT_07 => X"088C0060242183060CF118011281B00000220010400020002081A00082100001",
INIT_08 => X"40000400014812466427040098C000622AAAA43E3060C158AC97F0356BDBFBD0",
INIT_09 => X"00026C000559102400200281400469000008B0800000901080004004308B4340",
INIT_0A => X"045413002200000000400408200000201041000208000040020820034200005C",
INIT_0B => X"41E11C008089540000420100101088400000808404004000000020A000100414",
INIT_0C => X"18C191AC191A4191A4191AC191AC191A4191A00C8560C8D08400000609010100",
INIT_0D => X"0E08A20BC417C16004C0B8382210904018000080100100012200000064064019",
INIT_0E => X"0E0615C96000000010200000802100022008100408020401020040100142200E",
INIT_0F => X"C06100000021E300B000000781E00140018000000781E00140018000002430E3",
INIT_10 => X"68C381C00000024E0000000781E00140018000000781E0014001908400005E11",
INIT_11 => X"088400003C30F00C000000155800D00000003E21C0700000000F001180000004",
INIT_12 => X"4000260640900004A400081401A0000004041218503E40300600000048043180",
INIT_13 => X"00009A0001208C30800025200003D807E0000000007252016000904618400013",
INIT_14 => X"480160000F00C0E06100000012D2005100409520381C00000005920004C0C812",
INIT_15 => X"0004025000120850B8180625400400000010711200510004B414780400000055",
INIT_16 => X"1004010040002002080000000804000A0000000011A000100208C008611430A0",
INIT_17 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_18 => X"0401004010040100401004010040100401004010040100401004010040100401",
INIT_19 => X"5800050008000000000000000001004010040100401004010040100401004010",
INIT_1A => X"1451451451564090C69606492492C09A8C205148D757DF8A94102E0001063A29",
INIT_1B => X"BADD6EB75BADD6EB75BADD555555555555555555555555555555555555555145",
INIT_1C => X"FFE0000174BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974",
INIT_1D => X"F5D2AAAB555555400000000000000000000000000000000000000000000303FF",
INIT_1E => X"EFA2D17DEBAF7D1574BAAAFBFDFFFA2FFD74000855555FFFFFFC01FF087BE8BF",
INIT_1F => X"145557BFDEAA5500154AAAAAEBFF455D04175FF5D7FEAAAA002ABDEAA5D2EBFF",
INIT_20 => X"20BAAAD540145F7D5574BAAA8415400005540155F7D16AB45002EA8ABA005540",
INIT_21 => X"975EFF7AEBFF550055555FF55003DE00A2FFFFFEFAAD57DE00082AAAA00082A8",
INIT_22 => X"16AABAAAAEBFE10AAFBD7545F7D5554AA5D2ABDEBA082A821455D2EA8B455D2A",
INIT_23 => X"FFEABEFA2FBEAB455D7BD55FFFF84155FFFFFFFFF55AAAABFFFF5D556AB45A2D",
INIT_24 => X"000000000000175FFF7D140010FF84174BA552EBDEBA0004020AA5D04155FFAA",
INIT_25 => X"4BFBC51FF1471E8BEF55242FF47015A800000000000000000000000000000000",
INIT_26 => X"0B6AEBAEAA5D2EBDFFFBED17FEAAF7D5524AAA2F0BAF7FABDFC7E10005F525D7",
INIT_27 => X"55142A8708202FBD257F1C7550492490E17EAAA2AAB8F4515043DFC75575C700",
INIT_28 => X"03D1420AD000B420820AAE2DB6FB6DF7DFD5038ABA140A2D00554517DEBDB6FB",
INIT_29 => X"25555F8FFDE38087FC51C7F7AABFF55BC5B555C74B8A38E38085BE8B47A3A005",
INIT_2A => X"BA4AF555168B68FEDF6AB52AAABD21EF1C2FEA5FDEBDB505FA4920AFE10082E9",
INIT_2B => X"17AEB8BFF155552B6F5E8BFF1EFBFDBFF5FF1C00BF5D25475C7B7FEAFF45BEAA",
INIT_2C => X"00000000000000000000000000000151EAE3D542A004380124921D20BFFFA0AA",
INIT_2D => X"3D795000087BC01458AFBC11FF55516ABEFDD003EFE5093DC000000000000000",
INIT_2E => X"550434D555C53E0CE2AAA8742BA5D2ABDFFFF7D57DEAAFFD5420B2A2D37DB07A",
INIT_2F => X"F0851575FFAAFBDD5542B2EDD608897FD610D01151C610592A974BAFBAC28B55",
INIT_30 => X"100F3D68FFFAABAC20EF04003FE102400144ABAAFFF7DE772FDD56588042F72E",
INIT_31 => X"4EA0006BFE007E2E8315DD02F6A81A239501755F504BDF557D79431FD006EABA",
INIT_32 => X"03158517BD745AEAEA8FAF0C55EAF57FF957CAAA7FABF7DFD0C6A7DFFFA07FC0",
INIT_33 => X"964A92B403EE18D5408A6F2AFADF6900FFFF68BEFDFFB4B1FE5551141E78A028",
INIT_34 => X"0000000000000000000000000000000000000000000000165BAFBD542000D382",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000400000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0812",
INIT_01 => X"2145A00A1079284D04A044A54E504368404000720885800802000006ECD10200",
INIT_02 => X"5C010800020408040C415854AA055254090541A111000A104A00000009083510",
INIT_03 => X"0C1000100C0000D40526480250149120031500A0218808002440804288890550",
INIT_04 => X"8840C28120051400582012021808040409C0B26850488419444010C10A024A49",
INIT_05 => X"488510910548012025C0C0000300086854B141042252142042A048D090006372",
INIT_06 => X"948037480159A403109848000428AA8282102040449090D520085224410AA420",
INIT_07 => X"01020402242000408468112010810C055200022025A83AA3008882004A001542",
INIT_08 => X"11491C154429220A2824640010A010020282843E0008124C0000211000008840",
INIT_09 => X"E280442C1411D020828A2B116824632885419240016001900AE01A2020066395",
INIT_0A => X"30105108880684145002021012D40D718241108815380200900160AE42CE2818",
INIT_0B => X"53419F10308D100054AA080092112C100B400880454058E80B94080C49318000",
INIT_0C => X"D0090D0090D2890D0890D2890D0890D2090D0048610486808403A384880B8981",
INIT_0D => X"8202043800000620500403080A919000B8AD0304144008111A00582043243050",
INIT_0E => X"9835300002AA40AA902408200010002021060C810241832241280C81A0984020",
INIT_0F => X"100000000080A0000140000002000140200A8000000200014020100290E469C6",
INIT_10 => X"00100000000003400A8000000200014020094000000200014020087000000000",
INIT_11 => X"014200000004000000000081400004C00000000020000000008C000010A00000",
INIT_12 => X"0510000000000006800001880004008400800000000020000000000048100000",
INIT_13 => X"0000D0260000000000003409280000000000000040025000030000000000001A",
INIT_14 => X"400002A0000000000000000042900000A100000000000000008012A200000000",
INIT_15 => X"000000004420300000000000000000000010C010000098000000000000000105",
INIT_16 => X"00802208036408C0820010004D36A222120090554000E40080000000088000A0",
INIT_17 => X"8802008020080200822088220882208802008020080200822088220882208802",
INIT_18 => X"8320883200812008120081208832088320883200812008120082208822088220",
INIT_19 => X"E88051029FC0FC0FC1F81F81F820883208832088320081200812008120883208",
INIT_1A => X"08208208208C13A4301040B2CB2CBAC838B6C0080271AE180616A851158E2863",
INIT_1B => X"944A25128944A25128944A082082082082082082082082082082082082082082",
INIT_1C => X"FFE381F928944A25128944A25128944A25128944A25128944A25128944A25128",
INIT_1D => X"A550002000AA800000000000000000000000000000000000000000000003C200",
INIT_1E => X"BAFFAE801FF087BE8BFF5D7BEAA1055042AA105555421EFFFD568AAA002EBFEB",
INIT_1F => X"FFFA2D57DE10557BE8ABAF7AAA8BEFAAAE975FFA2D5555450851574000851554",
INIT_20 => X"5555F7D568ABAF7D5574BA552EA8AAA5D2EBFFFFA2D1554BAF7D17FEBAAAFFFD",
INIT_21 => X"EAAAA552AAAAAAAAAABFF455D04175FFFFD5574AAAAAA974BA082EA8BEFAAD55",
INIT_22 => X"FEAA000055401555D7BFFE10085557410F7AA97410087BD55FF087FEAA10A2FF",
INIT_23 => X"0017400550402155A2803FE005D7FE8B45F7FBFDE00085540155F7D56AA00007",
INIT_24 => X"00000000000017400082AAAA00082A820BAAAD540145F7D557410AA8428A1055",
INIT_25 => X"4BD16FAAA002ABFEAA550E82000E28A800000000000000000000000000000000",
INIT_26 => X"FEAFBD2410005F57482E3AA801FF1471E8BEF5574AFA00010ABFA38555F401D7",
INIT_27 => X"AAF7D5524AAA2F1FAF7FABFBFF400417FEF082F7AAA8BEFE2AA955EFA2DB5757",
INIT_28 => X"492082EADBFFBEDB55555E3DF6DA82F7DF520385D2FE80AA5D2EBDFD7BED1574",
INIT_29 => X"21C7005B6FB47F7A438E925D24ADAAAB6AAB8F455784155C75575C7000B6AE95",
INIT_2A => X"4717DEBDB6FA3D0075EDA800051C05571474024A81C5557578EBA087400007FC",
INIT_2B => X"FFDE381D716FA15550015428E10A001FFB40038F68F7F578F7FFEF568E280855",
INIT_2C => X"000000000000000000000000000001043D1420AD000B420820AAE2DB4716DF7D",
INIT_2D => X"828FDEBA5D7BC015582D57DEAA002ABDEAA552A80010AAA88000000000000000",
INIT_2E => X"AAAE955EFAAFBC15F5A3D7D6800087BD5410AAAA801FF55556ABEF5D517EEE00",
INIT_2F => X"A5D2ABDF55F7D575EAAFFD50A2B2A3D169B07A3D7BFE10597BFDE00AEAC28BFF",
INIT_30 => X"555A53C00B2A2AA02000082ABDFEFFFFBC1154AAFFFFE107FF9D72A20842080B",
INIT_31 => X"4EAA28015400547FC315D00797CF4780286A2105D2A3FEBAFFAC28B555504145",
INIT_32 => X"99ADABD5A8AAA0051575FFA2FFFDA02003FFDEAA8557D65550915544AA5D5157",
INIT_33 => X"144ABAAFFD75E7F2BDDD2B8016F9E2555500174AA282E20BFFFF842AAAAADD56",
INIT_34 => X"0000000000000000000000000000000000000000000000030EF04003FE102400",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000800000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380206",
INIT_01 => X"200C9A40408001683C0462C99E004B61404040028804A0080A000416A0990A0C",
INIT_02 => X"4809A900031800444461089866E331352180D468B8040E600C0081110B802CD0",
INIT_03 => X"6D0B61108C00014231A3080408C68420330066010A80881068A808401CC46330",
INIT_04 => X"482218066A09C03B348C1C1928DD5A4402211A68470944842640902107002D24",
INIT_05 => X"0583180353202020000144E50B44644B30A86D05014A0D224063095092100E34",
INIT_06 => X"54023740216934020303680A040066D98A182210085A50C02048288234629414",
INIT_07 => X"018C00220430814204E01C581291820CCA000E3226413990008C80205A00CCCC",
INIT_08 => X"4108747320081246252D5010184000220002A43E10294258E805E1156002D940",
INIT_09 => X"D0AA546AC41B112029A61D84424429AA1320B1010140C1350B48292020024180",
INIT_0A => X"000102022850A1CC0047071913208CE802430488082042008040F399606F4058",
INIT_0B => X"5141BE42B88840005268081412152900484201A814144D60888CAA2C48151020",
INIT_0C => X"1B49019490194901B4901B4901949019C901B64805E480CA94480506980125C4",
INIT_0D => X"5A01E2B1080602E00C54216800859000199C98800C8140A11A44423040240450",
INIT_0E => X"28A65300E6664599902600009821204A040C1C040C0205038300480801480208",
INIT_0F => X"000000000090000003202900000010002008A02900000010002008039666928B",
INIT_10 => X"00000000000801000A202900000010002009E0290000001000200A3800008000",
INIT_11 => X"036000008000000000000088000002D003008000000000000280100016200812",
INIT_12 => X"05B008088000008201021C880000488002810005000000000000040000100000",
INIT_13 => X"0010402B80412000000410199800040000000000408020000680209000000208",
INIT_14 => X"800012980040300000000000C020000C8300208800000000008200AE01011000",
INIT_15 => X"40A0000841003100010401000000000002008020000C38000200000000000120",
INIT_16 => X"10070300704028820801400068360424820185CCE0128010020000008088021C",
INIT_17 => X"0070100701007010050180501805018050180501805018070100701007010070",
INIT_18 => X"070140601007014060100701C040180501C040180501C0401807010070100701",
INIT_19 => X"4A81454A26AA555AAB554AAB5541C040180501C040180501C040180501406010",
INIT_1A => X"08208208209441D0B0000092492480AA2860607818F18E0C851428200B262C31",
INIT_1B => X"D4EA753A9D4EA753A9D4EA492492492492492492492492492492492492492082",
INIT_1C => X"FFD55E21A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8",
INIT_1D => X"FAA8000155080000000000000000000000000000000000000000000000000200",
INIT_1E => X"EFFFD568AAA002EBFEBA555142000AA802AA10F7D57FEAA557BE8B45A2D5555E",
INIT_1F => X"A10550402000AAD56AAAA557BC0155A280021EFA2FFE8B4555042AA105555421",
INIT_20 => X"0010AA842AAAAFFD542000FFD5574000851554AAFFAE801FF087BC01FF5D7FEA",
INIT_21 => X"7DE105551420BAF7AAA8BEFAAAE975FF005540145A2D157410AAD17DFFF5D040",
INIT_22 => X"03DEBAAAFFFDFEFAAD57DEAAF7AE975FF080428B455D7FFDEAA5D55574BA0051",
INIT_23 => X"AE800AA087BD5555552A821EF007FFFEAAAAD5554AA552EBFFFFA2D5554BAF78",
INIT_24 => X"000000000000020BA082EA8BEFAAD555555F7D568ABAF7D5574BA552E800BAAA",
INIT_25 => X"E975EAB6DBEDF575FFAA8E02155080E800000000000000000000000000000000",
INIT_26 => X"5EBAEADA38555F451D7EBD16FAAA002ABFEAA555E02000E28AA8A38EBD578E82",
INIT_27 => X"FF1471E8BEF5575EFA00012A87A38AAD56DA824975C217DAA84021FFAAF5EAB5",
INIT_28 => X"400BED57FFD7410E05038BE8E2DABAFFDB47412ABFE90410005F57482E3AA801",
INIT_29 => X"FEBA5D71D742A407FFFE00555F47082E3AAA8BEFA02A955EFA2DB5757FEAFBD2",
INIT_2A => X"BFFD7BED157482F7803AEAAA2F1FAF7FABFBEAE2AEBA4974871C043AB6D4975F",
INIT_2B => X"F7AE38497FC00BAB6A4850821C75D25C74920821D708757AE2AA3FFC04AA552E",
INIT_2C => X"0000000000000000000000000000007092082EADBFFBEDB55555E3DF6DA82F7D",
INIT_2D => X"AA8A8ABAAAD568A1020516ABFFFFFFD75FFAAAE8014500288000000000000000",
INIT_2E => X"AA80001FFAAD57EB55A2A8ABEBA5D7BD5545A2D57DEAA002EBDEAA557BC0010A",
INIT_2F => X"0087BD5410AAAA801FF5555629EF5C517EEE00828D74AAFBD57DE000057C21FF",
INIT_30 => X"EFA8FBC15E5A3D5D7400FFD57DF55082E974AAFFAABDEBA77FDD66A0ABBDC200",
INIT_31 => X"50555002ABFF54517EEB25D57C14100957FF6105D7BD5400AAAC28BFFAAAE955",
INIT_32 => X"FA42A3D7020BA5D2ABDF55F7D1554A8FFC42AA10A7D169F57ABD7FEEBAAA8415",
INIT_33 => X"C1154AAFFFFE10FFF9DF202096F014AAFF84154105555C215500000014558557",
INIT_34 => X"000000000000000000000000000000000000000000000015400082ABDFEFFFFB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000400000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204002",
INIT_01 => X"01039802000820491C00650E1E004340403008418984014902030906A8D10200",
INIT_02 => X"480108A000000000444048E41E80F00A41043118680002000800000009882390",
INIT_03 => X"06504110080000D0040608024010102026001260300000003080880208C000F0",
INIT_04 => X"9100E98268154C1AE0B01C160033B944028290285AE0DC38E02090E81C22E801",
INIT_05 => X"5C0F20B36F000109200044C401041C4CF21C48B433483C8242EAE1B0000074C4",
INIT_06 => X"100007000059800310086A1A0022E18780000140C9D9D0930000F228075A6071",
INIT_07 => X"00000000242000008461000810818403C100060064012E00048C82201800BC28",
INIT_08 => X"0048CC8F01090602202C0400008000002202243E400010480000211540008810",
INIT_09 => X"40E0DC1EB5191120C7BE7D152201612E80E891E0614041340838450020422111",
INIT_0A => X"30545DAD8C2E0982400603003200872003FB1408082840002044007846164E0A",
INIT_0B => X"43411D10118D1A04522E000498140C104B260DA0404003C08B6000AC01128000",
INIT_0C => X"C5010C3010C1010C3010C1010C1010C3010C140869808618850BE6305989AB80",
INIT_0D => X"100140302800108018840440028480001B8780800000003102045C3443043410",
INIT_0E => X"3080620481E0E18790012A001001026808000002020101028100200180080201",
INIT_0F => X"000000000010000005C0200000001000000C4020000000100000000380E4C308",
INIT_10 => X"00000000000800000D00200000001000000EC020000000100000086A20008000",
INIT_11 => X"012820008000000000000008000001B00100000000000000020000002AA00010",
INIT_12 => X"06D0000080000080000241D80000800442800001000000000000040000000000",
INIT_13 => X"0010003A00002000000400021800040000000000008010000B00001000000200",
INIT_14 => X"400005900000100000000000801000089000008000000000000200F800001000",
INIT_15 => X"00000000A500100000000100000000000200001000002E000200000000000020",
INIT_16 => X"000000C032700000022400444934240A8021B63C005108010004100098098010",
INIT_17 => X"C010080200401008000040300800004010000200C01000020040100802004030",
INIT_18 => X"02000000000100C0300400008000000300C0100C00000020080000C030000000",
INIT_19 => X"20240142325930C9A6CB261934C000200801004030040200800000030040100C",
INIT_1A => X"14514514514E98264686668A28A260521CC45140C700FC0A0002870980831A28",
INIT_1B => X"1A8D46A351A8D46A351A8D555555555555555555555555555555555555555145",
INIT_1C => X"FFD5E7D8341A0D068341A0D068341A0D068341A0D068341A0D068341A0D06834",
INIT_1D => X"A5D55420AA002A80000000000000000000000000000000000000000000000200",
INIT_1E => X"AA557BE8B45A2D5555EFAAD140155080000155FF843FFEFAA84001FF5D043FEA",
INIT_1F => X"000AA80001555D04174AA002A80010FFAE975FFAA80001EFA2AAAAA10F7D57FE",
INIT_20 => X"00BA5D51555EF002AA8BFFAAAAAAA105555421EFFFD568AAA002EBFEBA555542",
INIT_21 => X"82000AAD568AAA557BC0155A280021EFA2FFE8B45F78400145FF842AAAAA2AA8",
INIT_22 => X"BC01FF5D7FEAA105D0428B4500003DFEF080428B455D002AABA5D2AAAAAA5D2E",
INIT_23 => X"80154BAA2FBE8AAAF7AA821EFAAAAA8BEF552E820000851554AAFFAA801FF087",
INIT_24 => X"00000000000015410AAD17DFFF5D0400010AA842AAAAFFD542000FFD57DF55A2",
INIT_25 => X"A284051D755003DE92415F42092142E000000000000000000000000000000000",
INIT_26 => X"71C0A28A38EBD57DE824975EAB6DBEDF575FFAADE02155080E85145E3803FFEF",
INIT_27 => X"AA002ABFEAA555F42000E2AA851455D0A124BA002080010FFA4955C7BE8E021C",
INIT_28 => X"145F7802AABAA2A480092415B505D71424AABD7F68E2FA38555F451D7EBD16FA",
INIT_29 => X"AA824924AAA92550A07038BED56DA824975C217DAA84021FFAAF5EAB55EBAE82",
INIT_2A => X"55482E3AA801FF1471C01EF5575EFA00012ABFB6D080A3AFEF080A2FB45490E2",
INIT_2B => X"B6FA12ABAEBDF7DAA80104BAAAFFEAA00F7AE821D7B6A02FBC71D0E10010005F",
INIT_2C => X"0000000000000000000000000000010400BED57FFD7410E05038BE8E2DABAFFD",
INIT_2D => X"02897555A2803FFFFAA841754555043FE10087BC2000552C8000000000000000",
INIT_2E => X"FF8017545F7AE821455D2CAAABAAAD57DE1000516ABFFFFFBD75FFAAFFC01450",
INIT_2F => X"A5D7BD5545A2D57DEAA002EBDEAA557BC0010AAA895555042E820BA080400010",
INIT_30 => X"FFAAD57EB55A2A880155F7802AAAAAA8002010007FC0155D5022A955FFACBFEB",
INIT_31 => X"BEF002EBDF45542AAAA0008043CAB0552C97CAAFFD57DE000057C21FFAA80001",
INIT_32 => X"CFE55D2CC2000087BD5410AAAA801FF5555421EF58517EAB00028A9BEF002EAA",
INIT_33 => X"974AAFFAABDEBAF7FDDE6A0AA90FDFEFA280020BAA2FFEAA10FFAE82145F7803",
INIT_34 => X"000000000000000000000000000000000000000000000002000FFD57DF55082E",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000800000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A337A20E07C0C1E006",
INIT_01 => X"295FBC468000A04D5C6A60000C34C24841280A00084000C8C212892EEAD53235",
INIT_02 => X"C809AD5CB118E640A4D158F8011FF0002080000082C8C66609DB7DDDCB1F2036",
INIT_03 => X"250906263A4C904214A35C80085285720B20648A88800000B8E0F852A884500E",
INIT_04 => X"4005122126899100064D20001044429C78A43A2C4436CC87198A3916E0551A24",
INIT_05 => X"A370C14CA0E900004048402389CFE2F20F7D7A354CB5C208E51437F044948912",
INIT_06 => X"9B9407B9424F33468B096FCF452AE0505A185905CC2414D44437118630839B88",
INIT_07 => X"588C732074A68D5AB4EB180717FF513FC52691924098712CE481FDC201D43C1A",
INIT_08 => X"0016053F180A1286A4ED1BC18840C320000055FE91AA545CBA4DE1D17992D9BE",
INIT_09 => X"2D1A4D8105B734723041008100486100601EDE1DE46431138DFD404CB4022595",
INIT_0A => X"A131112C0D15C901B2122309204C28B67061E81A8920C8D3CF8014007902DA6B",
INIT_0B => X"AD5C3402488888E5126BA350B27C092E63D18C9C500577EEA33EF24C09B42464",
INIT_0C => X"096B80D6B80B6B80F6B8096B80F6B80B6B80D15C04B5C07AD50C94020D233107",
INIT_0D => X"8948020D829FA454104132252011E542387F810480C840C383751EF5606E0178",
INIT_0E => X"000200CA7FE0627FD25845E42151648F854480A042512028100A8C38280AA04C",
INIT_0F => X"D06101C55DE5E3E3C017E37FC3E0017C3F8817E37FC3E0017C3F900040241001",
INIT_10 => X"6CD381C0118797FE0817EA7FC3E0017C3F8817EA7FC3E0017C3F9900DFFFDE15",
INIT_11 => X"F800DFFFBE34F00C0270F3F55F1F8007FDBEBE25E0700463E1FF2C7E014FF7BE",
INIT_12 => X"C5DEF64EC090626FE40140459759173BBD6EF37D523E6030061341F07FD571F8",
INIT_13 => X"0C4DFE2A6FE2AC3082637F281BFFFC07E00007E07F7253D38337D1D6184131BF",
INIT_14 => X"4F4F8397FFA0F0E06101C53E76D3D3E884FDDDA8381C0098E5FD92BBDFC8D812",
INIT_15 => X"19074FA36FDF58DBF81C072540049707E0FEF313D3E03BFFF61478040570EFD5",
INIT_16 => X"8CA02ACA00C50850182309444D248204201040FC190054A2110B8ACC483204A1",
INIT_17 => X"0A128CA0284A2280A1288A128CA2284A0288A1288A3284A228CA0288A1280A32",
INIT_18 => X"A228CA0284A3280A3288A1288A3280A2284A028CA2284A2284A028CA0280A328",
INIT_19 => X"F6A1850E1892596D34924B2DA6A84A2284A1288A1280A3280A1288A0284A2284",
INIT_1A => X"7DF7DF7DF7CBFBFE7EFEEE79E79EFAF3F51EB769CFEF73B6FFE74FC2400DB6DB",
INIT_1B => X"EEF77BBDDEEF77BBDDEEF77DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF",
INIT_1C => X"FFC27F6BDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDD",
INIT_1D => X"55D2E955FFF7FFC0000000000000000000000000000000000000000000000200",
INIT_1E => X"EFAA84001FF5D043FEAA5D04020AA002AAAABA555140155087FFFFEF00042AB5",
INIT_1F => X"1550800001FF5D00001555D2E975FF5D5568B555D7BD5545FFD540155FF843FF",
INIT_20 => X"FF45A2FFC0000AAAE974AAFFFFEAA10F7D57FEAA557BE8B45A2D5555EFAAD540",
INIT_21 => X"401555D04174AA002A80010FFAE975FFAA80001EF002AAAABAF7D168A10A2D17",
INIT_22 => X"EBFEBA555542000A28028BFFF7803DF55FFAEBFE005D2EAAB45557BD55555555",
INIT_23 => X"517DF55082E974BA087FE8B55552E955EF5D7FEAA105555421EFFFD568AAA002",
INIT_24 => X"00000000000000145FF842AAAAA2AA800BA5D51555EF002AA8BFFAAAA820AA5D",
INIT_25 => X"007FFFFFF1C042FB7D492A955C7F7FBC00000000000000000000000000000000",
INIT_26 => X"5E3DB45145E3803AFEFA284051D755003DE92410F42092142E28ABA5D5B4516D",
INIT_27 => X"6DBEDF575FFAADF42155082E851C75D0E02145492E955C75D5F6DB55497BD554",
INIT_28 => X"ABAF7D16DA28A2DB7AF7DB6FBC7028A2AA95492FFFFE8A38EBD57DE824975EAB",
INIT_29 => X"FB45557BD5555415F45145490A124BA002080010FFA4955C7BE8E021C71C0A2D",
INIT_2A => X"451D7EBD16FAAA002ABFEAA555F42000E2AAA8BEFE3843AF55E3AABFE105520A",
INIT_2B => X"4821D7F68E07082495B7FF7D082E954AA087FEDB7D5D2A155D7157BEFA38555F",
INIT_2C => X"0000000000000000000000000000002145F7802AABAA2A480092415B505D7142",
INIT_2D => X"52CAAAAA5D7FD75EF087BFDFEF5D003DFEF002E95555F7FDC000000000000000",
INIT_2E => X"5D7BFDF45007FD7555A2F9D5555A2802ABFFAA841754555043FE10082A820005",
INIT_2F => X"AAAD57DE1000516ABFFFFFBD75FFAAFFC0145002895545552E80145002E95545",
INIT_30 => X"45F7AE821455D2CBFEAAFFD17FEAAAAFFEABFFF7FFD54BAA2AA95410F7FDEAAB",
INIT_31 => X"B45AAAABFE0009043FF555D7BD55550879D5555002E820BA080400010FF80175",
INIT_32 => X"75455D7DFFEBA5D7BD5545A2D57DEAA002EBDEAA557BC0000AAA8A8BEFA28028",
INIT_33 => X"02010007FC0155550222955FFAC97400087FFFFFF002E954AA087BFFFFF5D2E9",
INIT_34 => X"000000000000000000000000000000000000000000000000155F7802AAAAAA80",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000003000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B0061A258A2840112C03002C180004003220200403302301C0381A0086",
INIT_01 => X"860041C83839484C00A100000052024841000000090800090210010000510204",
INIT_02 => X"080108200C1000004464080400C0080100000000010432400800800009882050",
INIT_03 => X"040001008C2340D0800208624200002183800584488000103080010C08C10000",
INIT_04 => X"00101610A029B08400044800000000040008102A040810040400900500001800",
INIT_05 => X"02800000400C830934E4A0002900404400820000000A00824004084011200A00",
INIT_06 => X"14C8874C884D0C024608680210C11F8010122100880802800308010000829400",
INIT_07 => X"060800002430200004611000508184803A0900224000200008818028C04883E1",
INIT_08 => X"4041FE80E009024260240010608000000000043E040000488000201400008810",
INIT_09 => X"0002447E041B112020208010404029006FE0B081003204502000002068621191",
INIT_0A => X"35E5148B0D916BBE39049191200000200441048108000220002FC5FA60000148",
INIT_0B => X"5358BF12E88D1000022808801A112D1443142A815440600083FE9AA300100281",
INIT_0C => X"C1416C1416C5416C5416C3416C3416C7416C500B60A0B60AD40E34104C093904",
INIT_0D => X"8C03403C440C054048850A300A8480009A0020865AE4ECB11B441A105B05B016",
INIT_0E => X"00000031001E4800022100321489214001A742D3A368D1B4686D100234B44242",
INIT_0F => X"00000000000AB800302008000000014000602008000000014000674000260000",
INIT_10 => X"0000000000000241E020010000000140006020010000000140006A8400000000",
INIT_11 => X"028400000000000000000003C00052000200000000000000000CD00184000800",
INIT_12 => X"30000800000000049A48184000A0400000010000000000000000000048028C00",
INIT_13 => X"0000918480010000000024C9E000000000000000000FF0006440200000000012",
INIT_14 => X"C000602800400000000000000BB000112B0020000000000000007E0000010000",
INIT_15 => X"02A0005000202500010000000000000000104CF000198000000000000000000F",
INIT_16 => X"4AD2B46D180684E8402440044C24A30819020603E0A20640C8400010218432A0",
INIT_17 => X"2D1B4ED3B4AD0B42D1B4ED2B42D0B46D1B4ED2B42D1B46D3B4AD2B42D1B46D2B",
INIT_18 => X"D1B42D0B46D2B4AD1B46D0B4AD3B4ED0B46D1B4AD2B4ED1B42D0B4ED3B4ED0B4",
INIT_19 => X"F8840000331C618E38E38C31C7346D3B4AD3B46D0B42D3B4ED2B42D1B42D2B4E",
INIT_1A => X"1C71C71C71CEDBB676F66EFBEFBEFAF99CFEF179CFF1FE1E9F52AFF9BFAFBE7B",
INIT_1B => X"FE7F3F9FCFE7F3F9FCFE7F1C71C71C71C71C71C71C71C71C71C71C71C71C71C7",
INIT_1C => X"FFE43591FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"05D2EBDF55557FC0000000000000000000000000000000000000000000030200",
INIT_1E => X"55087FFFFEF00042AB555D2E955FFF7FFC21EFF7D17DEAA5D2AAAAAA5D557DE1",
INIT_1F => X"0AA002A82145555542010FF803DEAA5D5568BEF5D042AA10A2AAAAABA5551401",
INIT_20 => X"20BA00557DF455D7BFFEAA555540155FF843FFEFAA84001FF5D043FEAA5D0002",
INIT_21 => X"001FF5D00001555D2E975FF5D5568B555D7BD5545FFD568AAA5D00154AAAAD14",
INIT_22 => X"5555EFAAD540155080000000F7843FF55007FFDEAAA284020BAAAD168BFF0800",
INIT_23 => X"51401EFF7842AA00FF8417545AAAEBFE10FFFFEAA10F7D57FEAA557BE8B45A2D",
INIT_24 => X"0000000000002AABAF7D168A10A2D17FF45A2FFC0000AAAE974AAFFFFC21EF55",
INIT_25 => X"5520ADA92495B7AE10412EBFF45497FC00000000000000000000000000000000",
INIT_26 => X"0AAAAA8ABA5D5B4516D007FFFFFF1C042FB7D492A955C7F7FBC71EFFFD57FE82",
INIT_27 => X"D755003DE92410E02092140E0716D415F47000F78A3DE92415F6ABD7490A28A1",
INIT_28 => X"A92550A104AABED1470AA005F78F7D497FFFE925D5B45145E3803AFEFA284051",
INIT_29 => X"20BAA2DB68BC7140E051C75D0E02145492E955C75D5F6DB55497BD5545E3DB6A",
INIT_2A => X"7DE824975EAB6DBEDF575FFAADF42155082E87038FF8038F6D1C7BF8EAAAA800",
INIT_2B => X"A95492FFFFC71EF415F471C7FF8428A00E38412545AAAE3FE10A3FBE8A38EBD5",
INIT_2C => X"000000000000000000000000000002DABAF7D16DA28A2DB7AF7DB6FBC7028A2A",
INIT_2D => X"7FDD55EFF7D57DE005D003DE00007FEAA10002ABFF450079C000000000000000",
INIT_2E => X"087BE8B45082EAAA10A2A8AAAAA5D7FD75EF087BFDFEF5D003DFEF002E95555F",
INIT_2F => X"5A2802ABFFAA841754555043FE10082A82000552C955FF007BD5410FFAABFE00",
INIT_30 => X"45007FD7555A2F9EAA005D2A820AAF7D5574AA087BEABEF007FFDE00557DD555",
INIT_31 => X"BFF557BE8ABAA284020BAA2FBEAB55552C95545552E80145002E955455D7BFDF",
INIT_32 => X"FE10A2F9EAABAAAD57DE1000516ABFFFFFBD75FFAAFFC01450028974BAFF842A",
INIT_33 => X"EABFFF7FFD54BAA2AA95410F7FDD55EF007BD5555F7802AA10AA8000145AAAEB",
INIT_34 => X"00000000000000000000000000000000000000000000003FEAAFFD17FEAAAAFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000002400000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10800B0048201002842002C02450018800002300500030B313300C418992002",
INIT_01 => X"A34009C23838684D1C20E0000E11426840000000080000080200080000110200",
INIT_02 => X"4801082048100000446558040080000041000000000622400800000009000010",
INIT_03 => X"040001818CA144D0842248424210812103000480088000003080014688800000",
INIT_04 => X"000012002041900000048000000000040088322944200C850001940400301800",
INIT_05 => X"0200000040084000284000204104004402000025000800065004207030320800",
INIT_06 => X"108017080149000246086A2A1468004012120004440812D40120008200829001",
INIT_07 => X"2408000024302040846810005281848003494020400031240C8C8218E06A0009",
INIT_08 => X"4040050001090242602C0418408000000000243E0408104C8000201540008810",
INIT_09 => X"00024401041B132820000001424069004000B204636009104A0101226A422104",
INIT_0A => X"80049800A0281400300B0210200008B206639389480046240068180262000048",
INIT_0B => X"41401C1081811C44D22A18841616004118004482040448011800004D49340082",
INIT_0C => X"00192001920019200192041920419204192060C9010C90100008040008012101",
INIT_0D => X"48A000880144434A001001228000803198003604004048294008C40C483480D2",
INIT_0E => X"0000002160006000100000200811020805000480004000220108000060000800",
INIT_0F => X"09864038A2881210382000000001E003E0582000000001E003E0422834240000",
INIT_10 => X"0000160700706901982000000001E003E0582000000001E003E04E8400000000",
INIT_11 => X"0684000000000330C00F0C8210807200000000000581C01C1C809201C4000000",
INIT_12 => X"29D000000C2419121028C00020A2400000000000080082C180603A0E003A0904",
INIT_13 => X"8322414E800000432118908DF8000000061E001FC00C10207740000021908C48",
INIT_14 => X"40806BB800000009864038C14810201BAB000000026130071A80613A00000184",
INIT_15 => X"840080546520350000600812058100F81C018890201BBA0000008239020F1108",
INIT_16 => X"04812208033400C0022140404D268624B210040004A08400000044222900320C",
INIT_17 => X"0832048120481204822008020080204832048120480200802008020081204812",
INIT_18 => X"802008020C812048020080200812048120080200802048120483200802008020",
INIT_19 => X"0221054A2C208200010410400020880200812048120C80200802008120C81200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFD3B3D800000000000000000000000000000000000000000000000000000000",
INIT_1D => X"5AA8017410555540000000000000000000000000000000000000000000000200",
INIT_1E => X"AA5D2AAAAAA5D557DE105D2EBDF55557FFDE00557BEAABAA2AEAABEFF7801555",
INIT_1F => X"5FFF7FFD5555557BEABFFF7FBEAAAAAAD157555AA803FEBA5555421EFF7D17DE",
INIT_20 => X"DFEFAA80000BAAAAA820BAA2802AABA555140155087FFFFEF00042AB555D2E95",
INIT_21 => X"02145555542010FF803DEAA5D5568BEF5D042AA10A2AA955EFF7FFD5400F7FFF",
INIT_22 => X"43FEAA5D00020AA002ABDEBA5D7FE8A000004154BAF780001EFAAAAA8B450000",
INIT_23 => X"2AAABFF5551421FFAAD157545AAD5555EF557FC0155FF843FFEFAA84001FF5D0",
INIT_24 => X"00000000000028AAA5D00154AAAAD1420BA00557DF455D7BFFEAA5555575455D",
INIT_25 => X"AAA0A8BC7EB8417555AA84104385D55400000000000000000000000000000000",
INIT_26 => X"A4155471EFFFD57FE825520ADA92495B7AE10412EBFF45497FFFE385D71E8AAA",
INIT_27 => X"FF1C042FB7D492A955C7F7FBD056D5D75EABC7FFF5EAAAABEDF5257DAA8438EB",
INIT_28 => X"5EFEBFFD2400EBFBFAFEFAA80070BAA2A0870BAAA8028ABA5D5B4516D007FFFF",
INIT_29 => X"01D7AAA0AFB6D1C040716D415F47000F78A3DE92415F6ABD7490A28A10AAAA92",
INIT_2A => X"3AFEFA284051D755003DE92410E02092140E3DE924171E8A281C0E10482F7840",
INIT_2B => X"FFFE925D5B525454124AFBC74955421EFA2DF5557DAAD5D05EF0175C5145E380",
INIT_2C => X"000000000000000000000000000002AA92550A104AABED1470AA005F78F7D497",
INIT_2D => X"079FFEAA5D5568ABAA2842AB55A28015545A284000BA5D534000000000000000",
INIT_2E => X"F7FBC01EFA2842AABA0857555EFF7D57DE005D003DE00007FEAA10002ABFF450",
INIT_2F => X"A5D7FD75EF087BFDFEF5D003DFEF002E95555F7FDC01EF55556AB55F7D56AABA",
INIT_30 => X"45082EAAA10A2A8801FFA2FFC2000A2FFEABFFAA84174BAAA80174AAAA862AAA",
INIT_31 => X"AAA552A80010F78000145AA843DFEF5D02155FF007BD5410FFAABFE00087BE8B",
INIT_32 => X"21FF085755555A2802ABFFAA841754555043FE10082A82000552CBFE10085168",
INIT_33 => X"574AA087BEABEF007FFDE00557DC014500003FF450051401FFA2FBD55EFAAD54",
INIT_34 => X"00000000000000000000000000000000000000000000002AA005D2A820AAF7D5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00000648E2840112C00000418000002700500030B3132000400812082",
INIT_01 => X"A14008420008204D042100000212026840000000180800080200090048510204",
INIT_02 => X"080108000090000004655C040080000051000000000402400800000009000010",
INIT_03 => X"00000100803008D0842240024210810003800584488000103080894288800000",
INIT_04 => X"00009610A028B084000440C0040000040088323244280C950400808500321800",
INIT_05 => X"42800080400C8A09306420202804400402800035200A00020204287001114A00",
INIT_06 => X"14C8864C8849880002486800142BFF001292214444081254002801A200821400",
INIT_07 => X"004800002430204084281000D281040001182020400031241C0D80000041BFE9",
INIT_08 => X"444005000108020220240010048000000000043E0408104C8000000100008810",
INIT_09 => X"0812040105191100200081130210ED104008A285617205D02A01010141225091",
INIT_0A => X"8004C8252291490039039390200008B20E230008280040088040100240008061",
INIT_0B => X"40013C128BC95C44522A00241204094008442681100448000800826F49240001",
INIT_0C => X"0408000080000800008000080000800008000440020400229548040008012125",
INIT_0D => X"401140BC4028430108150900408590109A00209642E46CA00240460400200440",
INIT_0E => X"080410010000200002210A320C89000005A142D0A16850B6294D100234201242",
INIT_0F => X"2F9EC00000800008100020003C1FE00020080020003C1FE00020044014260082",
INIT_10 => X"132C7E3F00000100080020003C1FE00020080020003C1FE000200880000081EA",
INIT_11 => X"0080000081CB0FF3C000008000201000010001DA1F8FC0000080110080000010",
INIT_12 => X"040000B0BE6C00020040580040200000001004832CC19FCF81E0000000100002",
INIT_13 => X"80004020000C31CF60001000000007F01FFE00004000300420000618E7B00008",
INIT_14 => X"C0102000000F151F9EC0000040300401000200D547E3F00000800080001617AD",
INIT_15 => X"02A020100000822406E1B95A3F83000000008030040100000BAB87FB00000100",
INIT_16 => X"46D1B66D1A368C68D26000544D26A504AB120400222206404840001101843000",
INIT_17 => X"2D1B46D1B46D1B46D1B46D1B46D1B42D0B42D0B42D0B42D0B42D0B42D1B46D1B",
INIT_18 => X"D1B46D1B42D0B42D0B42D0B42D1B46D1B46D1B46D1B42D0B42D0B42D0B42D0B4",
INIT_19 => X"20840442200000000000000000346D1B46D0B42D0B42D0B42D0B42D1B46D1B46",
INIT_1A => X"3CF3CF3CF3DBF91E66C6FAD96D965201F4C251414A87D78AF421448BE28F3AEB",
INIT_1B => X"3E1F0F87C3E1F0F87C3E1F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"FFD160B27C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C3E9F0FA7C",
INIT_1D => X"AFFFFC2000557FC0000000000000000000000000000000000000000000000200",
INIT_1E => X"BAA2AEAABEFF78015555AA80174105555420000000021EFAA843DE00F7803FEB",
INIT_1F => X"F55557FD54AAA2AA955FF00043DE005504175FF08514014555557DE00557BEAA",
INIT_20 => X"DF45FFD17DFFFFFD56AA00557FC21EFF7D17DEAA5D2AAAAAA5D557DE105D2EBD",
INIT_21 => X"55555557BEABFFF7FBEAAAAAAD157555AA803FEBA55556ABFFA280154BAFF803",
INIT_22 => X"42AB555D2E955FFF7FFD5410002AAAAAAA2D57DF450004154BA087BEAAAAF7D5",
INIT_23 => X"843DE1008556AA00A28028B55FFD1555EFA2802AABA555140155087FFFFEF000",
INIT_24 => X"000000000000155EFF7FFD5400F7FFFDFEFAA80000BAAAAA820BAA280000AAA2",
INIT_25 => X"A2803AE38FF843DEBAEBFFC20285D75C00000000000000000000000000000000",
INIT_26 => X"55D5F7FE385D71E8AAAAAA0A8BC7EB8417555AA84104385D5542038000A001C7",
INIT_27 => X"92495B7AE10412EBFF45497FD24BAA2AA955C708003FE285D00155FF00554515",
INIT_28 => X"BEFA28E124AAF7843AF7DEBDB78FFFE3DF6DA284175C71EFFFD57FE825520ADA",
INIT_29 => X"04920875EAA82F7DB5056D5D75EABC7FFF5EAAAABEDF5257DAA8438EBA415568",
INIT_2A => X"4516D007FFFFFF1C042FB7D492A955C7F7FBD54380020ADA82BED57DF4508041",
INIT_2B => X"0870BAAA80070BAA2803DE00005F68A10BE802DB55E3DB555FFF68028ABA5D5B",
INIT_2C => X"00000000000000000000000000000125EFEBFFD2400EBFBFAFEFAA80070BAA2A",
INIT_2D => X"D53420BA082E82155AA802AAAAFF803DEBAAAFBC20BA55514000000000000000",
INIT_2E => X"5D04175EF0855575455D7BFFEAA5D5568ABAA2842AB55A28015545A284000BA5",
INIT_2F => X"FF7D57DE005D003DE00007FEAA10002ABFF450079C20BAAAAE9754500043DEBA",
INIT_30 => X"EFA2842AABA085768BFFA2AE820AAFF802ABEFAAFFEABEFAAFFFDEAA0051555E",
INIT_31 => X"E10F7D17FF5500000001008516AA10FFFFC01EF55556AB55F7D56AABAF7FBC01",
INIT_32 => X"75EFF7842AAAA5D7FD75EF087BFDFEF5D003DFEF002E95555F7FDD74BA08043D",
INIT_33 => X"EABFFAA84174BAAA80174AAAA86174AAAA843DE00087FE8A00F7843FF45AAFFD",
INIT_34 => X"0000000000000000000000000000000000000000000000001FFA2FFC2000A2FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000001000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000002300500030B3132000400812006",
INIT_01 => X"A1400802000020490000000000000240413C0A61590001D90213C90008510204",
INIT_02 => X"680108200010000054655C040080000041000000010402400800800009082011",
INIT_03 => X"00040100800020D0842240124210810043800504488000103081894288800000",
INIT_04 => X"00001410A00AA084000400C0060000040088323044201C850020820400101880",
INIT_05 => X"0200020040048A09202420000C00410402000025000800020804207000100800",
INIT_06 => X"10488704884D080202086A0A3429004012120004DC08125400A0008300821000",
INIT_07 => X"000800002C30204084381000128104000100002040003164040D800000400009",
INIT_08 => X"0440050003080202202400100080000000000C3E0408104C8000102300008810",
INIT_09 => X"4810240104111104200080120210A5104000A204615201500801010000AA10C0",
INIT_0A => X"81F525A82804010009029290200008B202238008080240000040100242048025",
INIT_0B => X"00A1141002C91844522A0004120488000800028000044000080020AF09240010",
INIT_0C => X"0408104081000810408100081040810008104040800408208040000008010121",
INIT_0D => X"4201E0B4000803200C150108008490809A002192462424202200440404204041",
INIT_0E => X"0804100160006000120002120499020A04A14650A32851962965190014200240",
INIT_0F => X"000000000080A200100021000000014020080021000000014020000014260082",
INIT_10 => X"0000000000000340080028000000014020080028000000014020008000008000",
INIT_11 => X"008000008000000000000081500010000100800000000000008C100080000012",
INIT_12 => X"05D0000880000006800058000020000000000005000000000000000048100100",
INIT_13 => X"0000D02E8040200000003401F80004000000000040026000274000900000001A",
INIT_14 => X"800023B8000030000000000042A00009AB00008800000000008012BA01001000",
INIT_15 => X"00A000106520350000040100000000000010C0200009BA000200000000000105",
INIT_16 => X"465196651B328CA8D26540544924272EB91004002022024048400000098030A0",
INIT_17 => X"6509425094250942509425094250942509425094250942509425094251946519",
INIT_18 => X"5094250942509425094250942519465194651946519465194651946519465194",
INIT_19 => X"2A05404808000000000000000014651946519465194651946519465094250942",
INIT_1A => X"69A69A69A68945B080201C92410480ABD102E689999E91BCD151200C30AE1C71",
INIT_1B => X"341A0D068341A0D068341A28A28A28A28A28A28A28A28A28A28A28A28A28A69A",
INIT_1C => X"FFC5B52068349A4D068341A0D269341A0D269341A0D068349A4D068349A4D068",
INIT_1D => X"0F7D17FFFFAAAE800000000000000000000000000000000000000000000003FF",
INIT_1E => X"EFAA843DE00F7803FEBAFFFFC2000557FEABEFA2D1400AA5D2AAAA00F7FFEAA1",
INIT_1F => X"4105555421EFF78028BEF5D003DFEFF7FFE8ABAF7802ABEFAAAE820000000021",
INIT_20 => X"AB45557BC0155007FFDEBAAA843DE00557BEAABAA2AEAABEFF78015555AA8017",
INIT_21 => X"154AAA2AA955FF00043DE005504175FF0851401455555555EFA2FBC01FFF7AAA",
INIT_22 => X"57DE105D2EBDF55557FFDE00552A974AAA2843DEAA5D2A820BA000428AAAAA84",
INIT_23 => X"517FFEFAAAEBDF45FFAEA8ABAF7D1400BAAAAE821EFF7D17DEAA5D2AAAAAA5D5",
INIT_24 => X"0000000000002ABFFA280154BAFF803DF45FFD17DFFFFFD56AA00557FC201000",
INIT_25 => X"4120ADA38E3F1EFA28F7DF7DFD7A2A4800000000000000000000000000000000",
INIT_26 => X"7A2A482038000A001C7A2803AE38FF843DEBAEBFFC20285D75EFBC7A2DB40082",
INIT_27 => X"C7EB8417555AA84104385D55421C7FF8028BEF41003FFD7F7F1EDA82F78E2DBD",
INIT_28 => X"5C7A2FBC51EFEBA0A8B6D5571C716D1475FFEAAA28E3FE385D71E8AAAAAA0A8B",
INIT_29 => X"50AA1C0428ABAB68E124BAA2AA955C708003FE285D00155FF0055451555D5F57",
INIT_2A => X"7FE825520ADA92495B7AE10412EBFF45497FFFE105D2E97482AA8038EAA412E8",
INIT_2B => X"F6DA284175C001000557FFEFB6A0BFF55F7AEAAA82FFDF40092B6A4871EFFFD5",
INIT_2C => X"0000000000000000000000000000028BEFA28E124AAF7843AF7DEBDB78FFFE3D",
INIT_2D => X"5517DF55A2FBC201008003DEAAA2D57FEAAF7FBFDF45AA800000000000000000",
INIT_2E => X"FFD57FE00FFAABFF45AA80020BA082E82155AA802AAAAFF803DEBAAAFBC20BA5",
INIT_2F => X"A5D5568ABAA2842AB55A28015545A284000BA5D5340145F78028BFF08003DF45",
INIT_30 => X"EF0855575455D7BD5555A2FBD75FFA2842ABFF5555575FF55557FEAAA2AABFEA",
INIT_31 => X"400A2802AABA002A954AA5D0028ABAF7AA820BAAAAE9754500043DEBA5D04175",
INIT_32 => X"2010FF80155EFF7D57DE005D003DE00007FEAA10002ABFF450079FFE005D2A97",
INIT_33 => X"2ABEFAAFFEABEFAAFFFDEAA00514200008517DFEFFF803FF45FFAAA8A00F7FBC",
INIT_34 => X"000000000000000000000000000000000000000000000028BFFA2AE820AAFF80",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000002000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800020030000000033022000000180006",
INIT_01 => X"0000098218302849180060000C00424040000000080000080200090008510200",
INIT_02 => X"0801080200100000044008000080000041000000002002400800000009008010",
INIT_03 => X"0001000004000040000202000000000803006400088000003080040008C10000",
INIT_04 => X"0000100022008000000C08C00C00000400201830040000040000000400001820",
INIT_05 => X"0200000040000000248080210044000400000000000800000004000010000800",
INIT_06 => X"100007000049000202086A080000004010100000880800001000000030829000",
INIT_07 => X"000800002420000004201000128100000300002040003124040D802040400009",
INIT_08 => X"040005000108020220240020008000000000043E000000488000000100008811",
INIT_09 => X"0810040105111000202000024010A51040088080000000110000002000020084",
INIT_0A => X"040000000000010000040010200008B202230480080002000000100240008021",
INIT_0B => X"40003C020AC04400022808001000014000040088140000000000828000000820",
INIT_0C => X"0040004400044000040000400044000440000400002000221048840009012124",
INIT_0D => X"0002A00800000100440000000800800018002000008000800040022000000400",
INIT_0E => X"0804100100002000100002001001024800020001000080004000000800904000",
INIT_0F => X"000000000000A000102008000000014000082008000000014000000000240082",
INIT_10 => X"0000000000000240082001000000014000082001000000014000028000000000",
INIT_11 => X"028000000000000000000001400012000200000000000000000C100084000800",
INIT_12 => X"0000080000000004800000400020400000010000000000000000000048000000",
INIT_13 => X"0000900000010000000024080000000000000000000250002000200000000012",
INIT_14 => X"4000200000400000000000000290000100002000000000000000120000010000",
INIT_15 => X"0000001000000000010000000000000000104010000100000000000000000005",
INIT_16 => X"0000000001400080002100544924002A000004000020000080000000010032A0",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100400000000",
INIT_18 => X"0000000000000000000000000010040100401004010040100401004010040100",
INIT_19 => X"02A1410808000000000000000000000000000000000000000000000000000000",
INIT_1A => X"145145145146AB2A0CCC2A28A28A7AA0CDF0D1215281FC1A72E24C28E921AAA9",
INIT_1B => X"CA6532994CA6532994CA65145145145145145145145145145145145145145145",
INIT_1C => X"FFD9C63B95CA6532994CA6532B95CAE572994CA6532994CAE572B95CA6532994",
INIT_1D => X"FAAD1555FFF78400000000000000000000000000000000000000000000000200",
INIT_1E => X"AA5D2AAAA00F7FFEAA10F7D17FFFFAAAE801FF08557DF4555516AA00007BEABE",
INIT_1F => X"000557FC0010AAD57FF45A2D56AA0000043FFEFA2FFFDE1008556ABEFA2D1400",
INIT_20 => X"DEAA007FEAB45AAAE800AAF784020000000021EFAA843DE00F7803FEBAFFFFC2",
INIT_21 => X"421EFF78028BEF5D003DFEFF7FFE8ABAF7802ABEFAAAEA8BFF5D0415400F7FBF",
INIT_22 => X"015555AA80174105555401FF5D0415555557BFDFEF00517DE00A28028B450855",
INIT_23 => X"FFD7555AAD56AB45A2AE800AA5D7FFDEBAF7AEBDE00557BEAABAA2AEAABEFF78",
INIT_24 => X"000000000000155EFA2FBC01FFF7AAAAB45557BC0155007FFDEBAAA8417410AA",
INIT_25 => X"55556AA381C75EABEFBED1575C7E380000000000000000000000000000000000",
INIT_26 => X"81C516FBC7A2DB400824120ADA38E3F1EFA28F7DF7DFD7A2A4801EF085F7AF6D",
INIT_27 => X"38FF843DEBAEBFFC20285D75C0010AADF7AF6DB6D56FA3814003AFFFA2F1F8E3",
INIT_28 => X"BEF550412428F7F5FDE920875E8B45BEA0850BAE38002038000A001C7A2803AE",
INIT_29 => X"8E10AA802FB450851421C7FF8028BEF41003FFD7F7F1EDA82F78E2DBD7A2A4AD",
INIT_2A => X"E8AAAAAA0A8BC7EB8417555AA84104385D55401C75504125455575FAFD714557",
INIT_2B => X"5FFEAAA28E10438AAF5D2545BED56FB45BEA082082557BF8EBAF7AABFE385D71",
INIT_2C => X"00000000000000000000000000000175C7A2FBC51EFEBA0A8B6D5571C716D147",
INIT_2D => X"A80021FF007BE8BFF5D516AABA5D5568BEFF7D157555AA800000000000000000",
INIT_2E => X"5D002ABFFA2D16AAAA55517DF55A2FBC201008003DEAAA2D57FEAAF7FBFDF45A",
INIT_2F => X"A082E82155AA802AAAAFF803DEBAAAFBC20BA555140010AAFFE8BFFFFD17DEBA",
INIT_30 => X"00FFAABFF45AA803FFEF5500020BAFFD17DE10005568B55FF80154BAA280020B",
INIT_31 => X"1555D556AB555D5568A00AA843FF55085140145F78028BFF08003DF45FFD57FE",
INIT_32 => X"AAAAF7AABFEAA5D5568ABAA2842AB55A28015545A284000BA5D5342145550402",
INIT_33 => X"2ABFF5555575FF55557FEAAA2AA800AAAAD142155F7D57DF45FF8002010557FE",
INIT_34 => X"000000000000000000000000000000000000000000000015555A2FBD75FFA284",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000023FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B830084C1820E0000C36424840000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"000406A492E6E440842254D002108153422004800880000030C0315688C00006",
INIT_04 => X"00001201200090001205400000000094108C322644240C840008030440111800",
INIT_05 => X"222000444008010028404002A002009402400025080880000C04223000170900",
INIT_06 => X"12801628014B0B000A086CA6556800C012121004540816544522008200821100",
INIT_07 => X"1C08320054B624408428100094ADD080011721A04000316C140CA1A8A1F90019",
INIT_08 => X"00140500090B02C2E0EC04D1C08000000000647E858A104C920C81A5011088A6",
INIT_09 => X"40002481041F165820000101024061004004800567603592A801014C46426011",
INIT_0A => X"8404002020000101B0070310200008B60A23A51B28024CE24E40100260040004",
INIT_0B => X"2800340208811865D22BB384100E01090805A495100400050800E24D49A424C5",
INIT_0C => X"0C72A0872A0C72A0872A0C72A0C72A0872A0C595043950421400800009010104",
INIT_0D => X"4290A088812203360410110A400085539800210404C048CAC040464D28014405",
INIT_0E => X"0804101160006000101004A01811064B050204810240812241280D00200A0804",
INIT_0F => X"6D0141B0482A01AAEC3602330CD2A02952DC3502330CB4A0318B414000240082",
INIT_10 => X"5B4551630144C0155C3502330CD2A02952DC3602330CB4A0318B5600C587149B",
INIT_11 => X"FE04E587083B6A51005956308D1E8202C436375908AA840AD4513437640F1524",
INIT_12 => X"E020C67062F47B2872400044959BC42B1060F0D036B80B548523136C158878D8",
INIT_13 => X"8F0B27010A2699AAA3794392000D81852B0A050C224180062085134CD1719564",
INIT_14 => X"0AD57400C50500D94C8121713C02B555101C90705D71009604140C0418CE0C37",
INIT_15 => X"DC06A27C828E024D8C50965A40821568A06113801505010334AA73AA0666DAC2",
INIT_16 => X"04812048123408C0822040004C248604B2100400100084008001D0113920060C",
INIT_17 => X"4812048120481204812048120481204812048120481204812048120481204812",
INIT_18 => X"8020080200802008020080200812048120481204812048120481204812048120",
INIT_19 => X"00A0014200000000000000000020080200802008020080200802008020080200",
INIT_1A => X"4104104104140D220A4A380000002A80E900C4C1100830181621409C80210821",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000410",
INIT_1C => X"FFC1F83800000000000008040000000000000000000201000000000000000000",
INIT_1D => X"0F7842AA00002A80000000000000000000000000000000000000000000000200",
INIT_1E => X"4555516AA00007BEABEFAAD1555FFF784020AAF7D542155F7D1400AAF7FFFDE0",
INIT_1F => X"FFFAAAEA8ABAFFD17FEBAFFAA800AA007FFDFFFA28428A000000001FF08557DF",
INIT_20 => X"00AAF78028AAAFF84020AAFFFBEABEFA2D1400AA5D2AAAA00F7FFEAA10F7D17F",
INIT_21 => X"40010AAD57FF45A2D56AA0000043FFEFA2FFFDE1008556AB45555568A10A2FFC",
INIT_22 => X"03FEBAFFFFC2000557FC0155FFD1555FF0804000AA000428A10AAAA801EFFFD1",
INIT_23 => X"8428A10087FD7400552EBDFEFA2FBFFF550000020000000021EFAA843DE00F78",
INIT_24 => X"00000000000028BFF5D0415400F7FBFDEAA007FEAB45AAAE800AAF78428B45A2",
INIT_25 => X"E3DF450AAF7F1FDE38FF8A2DA101C2A800000000000000000000000000000000",
INIT_26 => X"01C0E001EF085F7AF6D55556AA381C75EABEFBED1575C7E380000BAF7DB4016D",
INIT_27 => X"38E3F1EFA28F7DF7DFD7A2A4AFABAFFDF7AE82F7AA870AA0071F8FFFBE842DA1",
INIT_28 => X"B455D5B68A28A2FFC20AAEB842DAAAE38A02082E3FBEFBC7A2DB400824120ADA",
INIT_29 => X"8A28AAA4801FFE3DF40010AADF7AF6DB6D56FA3814003AFFFA2F1F8E381C516D",
INIT_2A => X"001C7A2803AE38FF843DEBAEBFFC20285D75C2145F7DF525EF140A050AA1C002",
INIT_2B => X"0850BAE3802DB6DAA8A28A00007FD74284120BFFFFBEF1F8F7D080A02038000A",
INIT_2C => X"000000000000000000000000000002DBEF550412428F7F5FDE920875E8B45BEA",
INIT_2D => X"A80020BAFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE10552E8000000000000000",
INIT_2E => X"085568BEFF7803FE10552E821FF007BE8BFF5D516AABA5D5568BEFF7D157555A",
INIT_2F => X"5A2FBC201008003DEAAA2D57FEAAF7FBFDF45AA803FEBAFFFBEAA00F7AE974BA",
INIT_30 => X"FFA2D16AAAA55517DF55557FEAAAAA2FFC00AAAA803FEAAA2AA82000A2FFFDF5",
INIT_31 => X"1EF552E974BA550028ABAA280001FFAAFFC0010AAFFE8BFFFFD17DEBA5D002AB",
INIT_32 => X"ABFF082E820BA082E82155AA802AAAAFF803DEBAAAFBC20BA555142155F7FFC0",
INIT_33 => X"7DE10005568B55FF80154BAA2803FFFFA2AAAAA00007FD74BA08003DFFFFFD16",
INIT_34 => X"00000000000000000000000000000000000000000000003FFEF5500020BAFFD1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000002000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C048000C048400380000007026040000000080000088200002802153231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"210D050012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"0080100022408000060DE0000066630C70241827041000040800820480001AA4",
INIT_05 => X"0240000C400000003C808003E0C8001401000000040900020904004000070800",
INIT_06 => X"1800068000491300CF0969A421C0004018184000100804005784000130821200",
INIT_07 => X"7E8C53200CA4850224301807D1CB45900147E03040083124FC0CD0C8A1FF0019",
INIT_08 => X"0046050013081206A4A503A9E8C0812000001C7E11A24058B84D40E33992D98F",
INIT_09 => X"010004810491175C20000080000821004010C01086003C13E000004EDF020400",
INIT_0A => X"000000000000010000180018200408B27E234913E9000CFA09A8180248001000",
INIT_0B => X"ACA0141000800021826933E03662802B3001E09F000000023000000000000867",
INIT_0C => X"0832F0C32F0832F0832F0C32F0832F0832F0C197861978400000000208010100",
INIT_0D => X"05FA0201E7F3F01F40401C17E800C7F3380020000000006AE01180493C5BC1AF",
INIT_0E => X"000200F500002200004005002001408400000000000000000000053A4096F807",
INIT_0F => X"246FC1B17B2C53F2FC16691DB587201EDDF4162B1DB527201EDDC46070241001",
INIT_10 => X"2A67DF2A01D5CC9794162B1DB587201EDDF416691DB527201EDDD884272592D6",
INIT_11 => X"288007258E995D5A825DBA569F9FF02547068618CD3CC45B7863AE7EC00D4B12",
INIT_12 => X"F6208C6CCA5C33717461C045B5B182019473D19D7CCD856106F31A683621BDFC",
INIT_13 => X"866E2FB10A652CC8E3538BBA01624E51AA6C0469AC5493F5688532966471A9C5",
INIT_14 => X"4F9B740041E1F5759001B4AA1853E6D5144AA9C914C8608D2724A4C4118D992B",
INIT_15 => X"DE07EAD9825682D4A36C0B0B4B85112B2C4A05D3E6D5051893335EB0072AA85A",
INIT_16 => X"00000000008000000821000048260020000004001DC0800000010E7F70171401",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0100401004010040100401004000000000000000000000000000000000000000",
INIT_19 => X"2A21010808000000000000000000401004010040100401004010040100401004",
INIT_1A => X"4924924924890380800016A28A28802B10B83728C1111026C152A23010848658",
INIT_1B => X"6432190C86432190C86432082082082082082082082082082082082082082492",
INIT_1C => X"FFDE003AC964B2592C964B2592C964B2592C964B2592C964B2592C964B2592C9",
INIT_1D => X"5FFAA80155F78400000000000000000000000000000000000000000000000200",
INIT_1E => X"55F7D1400AAF7FFFDE00F7842AA00002AAAA10FF8002155F7FFC200008041755",
INIT_1F => X"5FFF7842AB55080000145557FE8AAA080000155F7FFFDEAA0000020AAF7D5421",
INIT_20 => X"2000FF80020AAA2AAAABFF002E801FF08557DF4555516AA00007BEABEFAAD155",
INIT_21 => X"A8ABAFFD17FEBAFFAA800AA007FFDFFFA28428A00000028B4555043DFFFFFAE8",
INIT_22 => X"FEAA10F7D17FFFFAAAE80000A284174AAFF8428AAAFF8415545AAFBD7545F7AA",
INIT_23 => X"00000105D55400AA082A82155F7FFFDEAA08556ABEFA2D1400AA5D2AAAA00F7F",
INIT_24 => X"0000000000002AB45555568A10A2FFC00AAF78028AAAFF84020AAFFFBC215508",
INIT_25 => X"E3F5C000014041256DEBA487145F784000000000000000000000000000000000",
INIT_26 => X"2080E000BAF7DB4016DE3DF450AAF7F1FDE38FF8A2DA101C2AAFA00EB8E0516D",
INIT_27 => X"381C75EABEFBED1575C7E3802FB551C0E0516D417FEDA921C000017DEBF5FDE9",
INIT_28 => X"B55410A3FFC7F7A087000FF80070BAAAAAADBD70820801EF085F7AF6D55556AA",
INIT_29 => X"556DA2FBD7545F7AAAFABAFFDF7AE82F7AA870AA0071F8FFFBE842DA101C0E2D",
INIT_2A => X"400824120ADA38E3F1EFA28F7DF7DFD7A2A480000BE8A17482F78A28A92E3841",
INIT_2B => X"A02082E3FBC217D1C0E0500041554508208208017DF7F5FDE9208556FBC7A2DB",
INIT_2C => X"000000000000000000000000000002DB455D5B68A28A2FFC20AAEB842DAAAE38",
INIT_2D => X"52EBDE00AAAE975FFAAD1420005504001FFAA8015545F7800000000000000000",
INIT_2E => X"5504001FFAAD17DE00082E820BAFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE105",
INIT_2F => X"F007BE8BFF5D516AABA5D5568BEFF7D157555AA803DF45552E975EF007FFFE00",
INIT_30 => X"EFF7803FE10552EBDF45002EBFF55FF8017410FF84154BAAAAABFF450000021F",
INIT_31 => X"400F7AEA8A10A284175FFAAFBD5555F7AEBFEBAFFFBEAA00F7AE974BA085568B",
INIT_32 => X"DE1008517DF55A2FBC201008003DEAAA2D57FEAAF7FBFDF45AA8002000FFAE95",
INIT_33 => X"C00AAAA803FEAAA2AA82000A2FFC21EF552A954100851554000004021FFFFD17",
INIT_34 => X"00000000000000000000000000000000000000000000003DF55557FEAAAAA2FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00010100926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"0004122122029100100C00001200009C40A83A2044360C84190BAC04E0101820",
INIT_05 => X"027000004009050064C8C00104C10184034010250089C00EB004327064B60900",
INIT_06 => X"1B9416B94149000402086D42142800C012125804440812541027008230821380",
INIT_07 => X"0008320014B02848A4A8100015C55500057801A04000712C040CB1F880600009",
INIT_08 => X"005005000908020220E40170008042000000557E048A144C800590010000882D",
INIT_09 => X"0100250104B5310020000100020821004016CC1C616401910801010100CA2040",
INIT_0A => X"800000000000010192072310200028B6022346080802C0074AC0100259001004",
INIT_0B => X"A8201410008088C5D2288004120E802908800488000500050800404D49A42EB0",
INIT_0C => X"0400000000040000000000000040000000000000020000000000000008010102",
INIT_0D => X"4A02008000000360401021280800E400B800610C844848200028448400000000",
INIT_0E => X"000000086000600040D045E4195104D5854284A14250A12A512A880828984008",
INIT_0F => X"85D480949E07A80948354B6E68982167061037496E6838216706206810240000",
INIT_10 => X"652138E510B456587037496E689821670610354B6E6838216706220431961CA9",
INIT_11 => X"C2043196186A91674011CE61403562274AA49CD594CF00039C7C414B6509DA22",
INIT_12 => X"8A2E6A983014780CC8604040424A5323845932E620295879818170304B2F5002",
INIT_13 => X"8F019451654B9104A328665603148895D44E0251142B42A3D8B2A5C882519432",
INIT_14 => X"0AC5DC06A6C6A465AA0091482382B17614F2202858EE300991415B45CD530602",
INIT_15 => X"4000052E08DC8047F17D1C7C3C02128E587D6A02B17605A130A4E8BF00225885",
INIT_16 => X"84A1284A123508508220808048240604B2100C00022084809000D000393722A1",
INIT_17 => X"4A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A12",
INIT_18 => X"A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A1284A128",
INIT_19 => X"F1228154000000000000000000284A1284A1284A1284A1284A1284A1284A1284",
INIT_1A => X"75D75D75D75FFAFEFEFEEEAAAAAAFBF3FC1FF77DDFE7EFBEFFE7CFC0044FBEFB",
INIT_1B => X"FAFD7EBF5FAFD7EBF5FAFD75D75D75D75D75D75D75D75D75D75D75D75D75D75D",
INIT_1C => X"FFC0003BF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5",
INIT_1D => X"F007FE8A00AAFBC0000000000000000000000000000000000000000000000200",
INIT_1E => X"55F7FFC2000080417555FFAA80155F7842AB55552E821FFFFD5555EF552ABDFE",
INIT_1F => X"A00002A821EF5D7BC21FFFFFBD55EFAAD1554BA00556AA00AAD16AA10FF80021",
INIT_20 => X"FF45A2AABFEBA082A975555D55420AAF7D542155F7D1400AAF7FFFDE00F7842A",
INIT_21 => X"EAB55080000145557FE8AAA080000155F7FFFDEAA00002AB45082A821EF5D557",
INIT_22 => X"BEABEFAAD1555FFF7842AABAA2FFE8BEF5D517FF455D554214500043DEBAAAFF",
INIT_23 => X"AABDF555D2E955EFA28428A10552EBFEAAAAD1401FF08557DF4555516AA00007",
INIT_24 => X"00000000000028B4555043DFFFFFAE82000FF80020AAA2AAAABFF002E80000AA",
INIT_25 => X"EBD5525C74124B8FC71C71EFA28AAF5C00000000000000000000000000000000",
INIT_26 => X"8AAD16FA00EB8E0516DE3F5C000014041256DEBA487145F78428B6D4120851FF",
INIT_27 => X"AAF7F1FDE38FF8A2DA101C2A871C74975C01FFEBF5D25EFA2D555482085F6FA2",
INIT_28 => X"B7D1C24851FF495F7FF55A2A0BFE921C2E9557D415B400BAF7DB4016DE3DF450",
INIT_29 => X"214508003FEAABEFFEFB551C0E0516D417FEDA921C000017DEBF5FDE92080E2A",
INIT_2A => X"7AF6D55556AA381C75EABEFBED1575C7E38028A82B6F1E8BFF495F78F7D49554",
INIT_2B => X"AADBD7082087000AAA4BFF7D5D20905C7AA842DA00492EBFEAABED1401EF085F",
INIT_2C => X"000000000000000000000000000002DB55410A3FFC7F7A087000FF80070BAAAA",
INIT_2D => X"78028BFF0004175EFA2D54214508042AB455D517DEBAA2D54000000000000000",
INIT_2E => X"AAD557410007BFDEAAA2D57DE00AAAE975FFAAD1420005504001FFAA8015545F",
INIT_2F => X"AFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE10552E975450051401EFA2D5421EF",
INIT_30 => X"FFAAD17DE00082EA8BFF5504175FF087BFFF45AA843FE005D2A955FF087BC20B",
INIT_31 => X"BFF087BEABEF00554215500003FEBAFFFBFDF45552E975EF007FFFE005504001",
INIT_32 => X"FEAAFFD5421FF007BE8BFF5D516AABA5D5568BEFF7D157555AA8028A00FFD16A",
INIT_33 => X"17410FF84154BAAAAABFF45000017410AA803DFEF550402155A2843FE00082AB",
INIT_34 => X"00000000000000000000000000000000000000000000003DF45002EBFF55FF80",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000033FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"000103A7A00904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000120122009000100C00000000000400A83A2044200C840000800400101820",
INIT_05 => X"020000004008010024C0C0010040000402000025000800020004207000100800",
INIT_06 => X"108016080149080002086807542800C012120004440812541020008230821000",
INIT_07 => X"4008120054B42850B42A100010ED1500010001A040003164040CF5E201400009",
INIT_08 => X"00400500090A020220A40A7000800000000014FE8508144C924080C100008801",
INIT_09 => X"0000040104111100200001000200210040008004616001910801010000422000",
INIT_0A => X"800000000000010190070310200008B202236D080802400002C0100240000000",
INIT_0B => X"0000141000800844522800041204000008000488000400000800004D49240820",
INIT_0C => X"0400004000000000000004000000000000004000000000000000000008010100",
INIT_0D => X"42020080000002204010010808008000B8002104044048200000440400000000",
INIT_0E => X"0000000000006000000000201811004005020481024081224128080820984000",
INIT_0F => X"CBA340480040A100A42008000161C140000420080001C1C14000032010240000",
INIT_10 => X"1A8A039600022260042001000161C140000420010001C1C140001604E8084341",
INIT_11 => X"1E04E8082580E2B8802201014800C220A21829A302F1C024010C001124020C8C",
INIT_12 => X"0024ACA60CA000048228404401004418012787124648157780120B8678C00080",
INIT_13 => X"00009001072D04730000241000CB1325E78E0186030240000083B60239800012",
INIT_14 => X"00001001EF6F4163C480481506800004000CFD55196CB012481812049495C194",
INIT_15 => X"40068248800108B8FB61A0401200845594965000000400568D0CFB7800550605",
INIT_16 => X"04812048123408408220000048240604B210040000008400800B0000090022A1",
INIT_17 => X"4812048120481204812048120481204812048120481204812048120481204812",
INIT_18 => X"8120481204812048120481204812048120481204812048120481204812048120",
INIT_19 => X"2820014000000000000000000020481204812048120481204812048120481204",
INIT_1A => X"3CF3CF3CF3CFFBBEEEEEFE79E79EFAABDDFAF369CB91FE1EF7D3AEBBDBAFBEFB",
INIT_1B => X"FE7F3F9FCFE7F3F9FCFE7F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"FFDFFFC1FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"AAAAEAAB45082E80000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFD5555EF552ABDFEF007FE8A00AAFBE8BEFA2D568ABA00003DF555555574A",
INIT_1F => X"155F78428AAA007FE8A1008002AABA555155400557BC2010557BEAB55552E821",
INIT_20 => X"FFFF082EBDEBAA2D1420105D002AA10FF8002155F7FFC2000080417555FFAA80",
INIT_21 => X"C21EF5D7BC21FFFFFBD55EFAAD1554BA00556AA00AAD140145AA8028ABA002EB",
INIT_22 => X"FFDE00F7842AA00002A80155A2AEA8A10080428A10FFAEBFFEF5D0428B45A2FF",
INIT_23 => X"5568A000000175FFF7D155545F7FBC0010FFAA820AAF7D542155F7D1400AAF7F",
INIT_24 => X"0000000000002AB45082A821EF5D557FF45A2AABFEBA082A975555D55400BA00",
INIT_25 => X"000E38F6D4155504AAA2AEAAB6D0024800000000000000000000000000000000",
INIT_26 => X"05D75E8B6D4120851FFEBD5525C74124B8FC71C71EFA28AAF5E8BFFB6D56DA82",
INIT_27 => X"0014041256DEBA487145F78428ABA147FEDA10080E2AAAA555552400417FC200",
INIT_28 => X"155BE8028A82002EB8FC70024BAEAAB6DB4202849042FA00EB8E0516DE3F5C00",
INIT_29 => X"DFD7550428B55A2F1C71C74975C01FFEBF5D25EFA2D555482085F6FA28AAD147",
INIT_2A => X"4016DE3DF450AAF7F1FDE38FF8A2DA101C2A80145B6AEA8A10080E2DA00F7A0B",
INIT_2B => X"E9557D415B400AA00556DA000004175FFE3D15757DE3F5C0038FFAA800BAF7DB",
INIT_2C => X"000000000000000000000000000002AB7D1C24851FF495F7FF55A2A0BFE921C2",
INIT_2D => X"2D568BEFFFD57FE10002AAABEF0051400AAA2AAAABFF08000000000000000000",
INIT_2E => X"5D5142000007BC20105D5568BFF0004175EFA2D54214508042AB455D517DEBAA",
INIT_2F => X"0AAAE975FFAAD1420005504001FFAA8015545F78028AAA557FFFE00082EAAAAA",
INIT_30 => X"10007BFDEAAA2D557555FF8028A00082EAAB45000028ABAFFFBC20AA08043DE0",
INIT_31 => X"A10002ABFE00F7803FF555D002AB55AAD1575450051401EFA2D5421EFAAD5574",
INIT_32 => X"20BAFFAE820BAFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE10552E82155FFAAA8",
INIT_33 => X"FFF45AA843FE005D2A955FF087BC20AA00517DE000804175EFAAD1555EFA2D14",
INIT_34 => X"000000000000000000000000000000000000000000000028BFF5504175FF087B",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000080000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"0001100024A0800000440000000000040088322044200C840000011400151800",
INIT_05 => X"A200014C4000000020000000000B8094020000254C8800000514203000108800",
INIT_06 => X"10000600004B0044020868021428004012120005540812540020008600831000",
INIT_07 => X"00086100043224489428100010811100010001A040003124040CAC6000400009",
INIT_08 => X"00160500090A0282A06400100080C300000005BE0488104C8000000100008800",
INIT_09 => X"00000581041110022000000002002100400080046140011008010100008A0400",
INIT_0A => X"800000000000010180060210200008B2022304080800400007C0100240000000",
INIT_0B => X"0004140000800844522800041004000008000080000400000800000D09240000",
INIT_0C => X"0400004000040000400000000000000000004000020000200000000008010100",
INIT_0D => X"4A00008000000260001001280000C400B0002000000000000000440400000000",
INIT_0E => X"0000000840006000000000001001004004000000000000020100000000000000",
INIT_0F => X"0000000000000000002021000000000000002021000000000000046000240000",
INIT_10 => X"0000000000000000002028000000000000002028000000000000020000008000",
INIT_11 => X"0200000080000000000000000000020001008000000000000000000004000012",
INIT_12 => X"0020000880000000006000400080C0000000000D081202800000000000000000",
INIT_13 => X"0000000100402000000000100000040200100000000000000080009000000000",
INIT_14 => X"0000100000003088014000000000000400000088221100000000000401001000",
INIT_15 => X"4000000800000000048407170500000000000000000400000200000000000000",
INIT_16 => X"00000000023000000220000048240404A010040000008000000000000000020C",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0020014000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000020000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFC0000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"555003DE10A2FBC0000000000000000000000000000000000000000000000200",
INIT_1E => X"BA00003DF555555574AAAAAEAAB45082EBFE000004020AA552E80000F7FBC214",
INIT_1F => X"A00AAFBFDEBA555568BEFA2FBE8A10F7802AA0055003FE10007BE8BEFA2D568A",
INIT_20 => X"55EFF78428BEFAAD17DF55AAAEAAB55552E821FFFFD5555EF552ABDFEF007FE8",
INIT_21 => X"28AAA007FE8A1008002AABA555155400557BC2010557BFFFEFA2FFC20005D2A9",
INIT_22 => X"417555FFAA80155F7843DF455D2AA8B45AAD57FF55A2FBC21FFA28415400FF80",
INIT_23 => X"514200055002AA00AA802AABA002E9740055516AA10FF8002155F7FFC2000080",
INIT_24 => X"00000000000000145AA8028ABA002EBFFFF082EBDEBAA2D1420105D003FFFF08",
INIT_25 => X"412A87010E3F5C0145410E3DE28B6FFC00000000000000000000000000000000",
INIT_26 => X"8147FE8BFFB6D56DA82000E38F6D4155504AAA2AEAAB6D0024B8E381C0A00092",
INIT_27 => X"C74124B8FC71C71EFA28AAF5F8EAA495F68BFFA2F1EFA38E38428A005D0038E2",
INIT_28 => X"FFFBEF5C0000492A955FFF78428BEFB6DB7DF45AAAEA8B6D4120851FFEBD5525",
INIT_29 => X"21EFAA8E10400E38E28ABA147FEDA10080E2AAAA555552400417FC20005D75F8",
INIT_2A => X"0516DE3F5C000014041256DEBA487145F7843FF7D4120A8B6DAAD17FF55B6F5C",
INIT_2B => X"B4202849043FFC7005F4501041002FA38A2842AA82142095428415F6FA00EB8E",
INIT_2C => X"0000000000000000000000000000007155BE8028A82002EB8FC70024BAEAAB6D",
INIT_2D => X"8002AAAA5D2A82000082E95400A2D542155002ABDEBAF7FBC000000000000000",
INIT_2E => X"A2802AA105D002AABA5D7BE8BEFFFD57FE10002AAABEF0051400AAA2AAAABFF0",
INIT_2F => X"F0004175EFA2D54214508042AB455D517DEBAA2D56AABA087BEABEFAAD57DEAA",
INIT_30 => X"00007BC20105D556ABFFF7D142010082A955EFFF8428BFFFFFBFDF55A2AEA8BF",
INIT_31 => X"BEFA2D57DF45F7D1401FFA2AA82000AAAAA8AAA557FFFE00082EAAAAA5D51420",
INIT_32 => X"54AA007BFDE00AAAE975FFAAD1420005504001FFAA8015545F7803FFEF08002A",
INIT_33 => X"AAB45000028ABAFFFBC20AA08043FF55087BD740000043DEAAA2842AA005D001",
INIT_34 => X"000000000000000000000000000000000000000000000017555FF8028A00082E",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000003000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"010108A802BB00080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"8BFA58800005C40A46240252145148B38248030356415A4E62B6FC660F287240",
INIT_05 => X"0F05EA11E570000D610000000710296E542B6E3A825C15FB30A643695BFC2D56",
INIT_06 => X"00000200021100C87570B08224C8AB52C0A8030140BCC0460050690A95C8383D",
INIT_07 => X"76F500240510A00205F0A407D0021A155378900002A002433A0AA00EE6E79564",
INIT_08 => X"00015995440C8327241440096A2800002828123D542910380004E03103624040",
INIT_09 => X"0010222D90409A05B2CB2CA400200209E5601044A24000000462A60018880100",
INIT_0A => X"300000000000259200140001A15000017F0051D0F837248C005514AC40C08205",
INIT_0B => X"395012004240014891801000495D40192D100000000005452D54000C09070003",
INIT_0C => X"6110001100011000110001100011000110001080008800080005202280801080",
INIT_0D => X"BB4000140A80A5C8000102ED0044008004AD324000000008003561180063DB4F",
INIT_0E => X"1400404912AA28AA890BA00000024800480000000000000200802151025062C0",
INIT_0F => X"6D0031F554E11C596A64003195933741477264003195555B418687E358360208",
INIT_10 => X"41CD50A499CF47DCB264003195933741597264003195555B4198843940076D29",
INIT_11 => X"043D400758486A556489347FE5F409CBC1362510695B6288743123C952518520",
INIT_12 => X"B1C74424EAE2992046EB70026486035600CEC45CBCA809654B48163CCC895E1E",
INIT_13 => X"C383298E3A242DEA151848302BFD6D522B10C7EC71F6C1DB071D1216E078C4C1",
INIT_14 => X"8B93D037DAAABC982BE22267A2E2E4F44AA1DC5E37400C9EE1B7B638E8849D23",
INIT_15 => X"86E6A2EE015998B28654565A003F0068E35352C1CAE48BFBF3A6C9B7B286B4DA",
INIT_16 => X"00000000009000040A8000452110A8442040D655602A102A0027E2C423202840",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"B020000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"28A28A28A28F4EF2FC3C34F3CF3C2AC31DF7A22A898D21B4C9838D30B6A7B451",
INIT_1B => X"F4FA3D3E8F4FA3D3E8F4FA68A68A68A68A68A68A68A68A68A68A68A68A68A28A",
INIT_1C => X"FFC00003E9F4FA7D3E9F47A3D1E8F47A3D1E8F47A3D3E9F4FA7D3E9F4FA7D3E9",
INIT_1D => X"AFF80001FF002A80000000000000000000000000000000000000000000000200",
INIT_1E => X"AA552E80000F7FBC214555003DE10A2FBC21FFFFFBFDF45A2D56AB45FFFFD54B",
INIT_1F => X"B45082E974BA5D7BFDF55A2FFFFE005D7BC0010002E954AA087FFFE000004020",
INIT_20 => X"7410FFD1555550000020BAAAFFE8BEFA2D568ABA00003DF555555574AAAAAEAA",
INIT_21 => X"BDEBA555568BEFA2FBE8A10F7802AA0055003FE10007BC0000082A9740055001",
INIT_22 => X"ABDFEF007FE8A00AAFBD55EFAAFBD74105504021FF5D2EAAABAFFFBD55FF002A",
INIT_23 => X"517DF45AAFFFFEAAFFAABFE10007FC00AA087FEAB55552E821FFFFD5555EF552",
INIT_24 => X"0000000000003FFEFA2FFC20005D2A955EFF78428BEFAAD17DF55AAAE820AA5D",
INIT_25 => X"AADB6FB6DFFFBD54AAE38E021FF0824800000000000000000000000000000000",
INIT_26 => X"A1C7FF8E381C0A00092412A87010E3F5C0145410E3DE28B6FFC21C7E3F1F8F55",
INIT_27 => X"6D4155504AAA2AEAAB6D002492482497BFDF45AAFFF8E385D7BC5000002E904B",
INIT_28 => X"010142E90428490015400FFDB555450804070BABEF5E8BFFB6D56DA82000E38F",
INIT_29 => X"DAAAFFF1D55FF002EB8EAA495F68BFFA2F1EFA38E38428A005D0038E28147FC2",
INIT_2A => X"851FFEBD5525C74124B8FC71C71EFA28AAF5D25D7B6F1D54384904021FF5D2AA",
INIT_2B => X"B7DF45AAAE820925D5B7DF45A2F1FDEAAEBAABDE001471C20921475E8B6D4120",
INIT_2C => X"0000000000000000000000000000038FFFBEF5C0000492A955FFF78428BEFB6D",
INIT_2D => X"7FBC2145AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF00000000000000000000",
INIT_2E => X"557FD7410082A800AA557BEAAAA5D2A82000082E95400A2D542155002ABDEBAF",
INIT_2F => X"FFFD57FE10002AAABEF0051400AAA2AAAABFF080000000087BFDF55A2FFE8AAA",
INIT_30 => X"105D002AABA5D7BC20005D2E800BA080417400F7FBD75450800174AAFFD168BE",
INIT_31 => X"4AA0800001EF5D2ABDEBAF7D1575EF082EAAABA087BEABEFAAD57DEAAA2802AA",
INIT_32 => X"0000555568BFF0004175EFA2D54214508042AB455D517DEBAA2D540155F7D155",
INIT_33 => X"955EFFF8428BFFFFFBFDF55A2AE82010557FFDF55A2D57FEAAAAAEBFE1055514",
INIT_34 => X"00000000000000000000000000000000000000000000002ABFFF7D142010082A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000001000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"294ADB4AFFCBF0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"DB7A40806FE4040840EBC563A0150A0926146FECB04196482236FC2005282AE1",
INIT_05 => X"0403DA0383200831C68206D7E6D0250834336D1E81500FDB306045255BFC2076",
INIT_06 => X"D0002200022D1C59E53558D3EBFC6701CBC303163670497AFF00291B3C0E2015",
INIT_07 => X"F81684248A38B022475DCA9BD00116E33CC3821774BB55F53BB42329AA3C0CEA",
INIT_08 => X"1660700CE0641527241060AD844E1C0088001223022D189A2800542219204903",
INIT_09 => X"B6D94C1C1C51DFF881861CBE0305A12A0321810217C01D34EDC98FFA1C8E0000",
INIT_0A => X"F1F1FD8F8FBDE40E001E000B3A5DAADAFDDA5DA79350DF70027CE86F047BEF19",
INIT_0B => X"2DD8141817C00319F8E853E64D73A08BFF00E9A7415606747E6610052CDEE97F",
INIT_0C => X"4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBCF4FBE7A7DE7A7800617112E46F05D0",
INIT_0D => X"BFF252D4CFEB69FF7A5F5AFFCCA787F7FE67C2180000006CE8A3F06ABD73DBCF",
INIT_0E => X"94BB02C9F99FD0678B87A0003000D8D02E00000000000000040025D3C21463D6",
INIT_0F => X"6D2BF232221ABD9CA854DFDD64A67D42C0F054DFDD64667D42C063E57A8F7B45",
INIT_10 => X"EFBB5AEDAA504801F054DFDD64A67D42C0F054DFDD64667D42C07237DFE5865F",
INIT_11 => X"3A33DFE58EAE7F5AB50D0806A9A2E0DFFF47DEDC496DA3181A0CC71440F9FBC3",
INIT_12 => X"7056E9C9C3FC95949AEFF556EF9C75E7DCF1EB1B6E6FCDC87CB35FC94B36AECF",
INIT_13 => X"92B29382AF5B6AAAE594A4C0DBFDAD94AA669809809FEFAF4157ADB55572CA52",
INIT_14 => X"BEBF41AE33F32ADD543430808BABAF50E1A5EB4BAEA45A250202FE0ADD39387F",
INIT_15 => X"E83FB669523E865D4B1293AB6B90BF2F0E30EDEFAFD0B3FBD72E9E90D20A003F",
INIT_16 => X"0000000002F840000BCE0B6F67B3F845E017C833F6AAC02B002A2EFF22D4073D",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"CC0C006000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"34D34D34D352324C3434C0EBAEBA21BBE5F04006013DB9880A5D25C3230B88A7",
INIT_1B => X"1A0D06A351A0D06A351A0D34D75D34D34D75D34D75D34D34D75D34D75D34D34D",
INIT_1C => X"FFC00002351A8D46A351A8D46A351A8D46A351A8D468341A0D068341A0D06834",
INIT_1D => X"0007BEAB55FFAA800000000000000000000000000000000000000000000003FF",
INIT_1E => X"45A2D56AB45FFFFD54BAFF80001FF002A821FFFFFFFFFFFFFFBFDFEFAAD14201",
INIT_1F => X"E10A2FBEAB45A28000010082A975EFA2D140145007BC21FF5D2A821FFFFFBFDF",
INIT_20 => X"54AA0855575FFAAD57FE005D7BFFE000004020AA552E80000F7FBC214555003D",
INIT_21 => X"974BA5D7BFDF55A2FFFFE005D7BC0010002E954AA087FD7400082E954AA08001",
INIT_22 => X"5574AAAAAEAAB45082EBFFFFF7D16AB45FFFFEABEF007BD74005555555EFF7AE",
INIT_23 => X"84154BA082E801FFAAFBC0155555568B45552EA8BEFA2D568ABA00003DF55555",
INIT_24 => X"00000000000000000082A97400550017410FFD1555550000020BAAAFFC0145AA",
INIT_25 => X"F7F1FAFD7A2D5400001C7BEDB7DEBA4800000000000000000000000000000000",
INIT_26 => X"F4124821C7E3F1F8F55AADB6FB6DFFFBD54AAE38E021FF0824851FFFFFFFFFEF",
INIT_27 => X"10E3F5C0145410E3DE28B6FFEFB45AA8E070281C20925FFBEDB451451C7BC01E",
INIT_28 => X"4280024924AA1404174AA0055505EFBEDB7AE385D7FF8E381C0A00092412A870",
INIT_29 => X"54005D5B575EFEBAE92482497BFDF45AAFFF8E385D7BC5000002E904BA1C7FD5",
INIT_2A => X"6DA82000E38F6D4155504AAA2AEAAB6D0024BFFD7FFDB6AB7DFFF5EDBC71C7BD",
INIT_2B => X"4070BABEF5C516DAA8A124921C20801FFB6F5C0145555B68B7D4124A8BFFB6D5",
INIT_2C => X"0000000000000000000000000000002010142E90428490015400FFDB55545080",
INIT_2D => X"000155FFF7FBFDFEFFFD568B45AAD5400005D7BFFFEFAA800000000000000000",
INIT_2E => X"FFFFD5545557BC21FF080002145AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF0",
INIT_2F => X"A5D2A82000082E95400A2D542155002ABDEBAF7FBFDF55A2AA974AA5D04001EF",
INIT_30 => X"10082A800AA557BD74BA0004000AA5500174AA0855421FFFFFBEAAAA5D7BEAAA",
INIT_31 => X"BFFF7D57FF455D7FD54105D7BD75FFAAAA80000087BFDF55A2FFE8AAA557FD74",
INIT_32 => X"8BEF000028BEFFFD57FE10002AAABEF0051400AAA2AAAABFF08003FF55F7FFEA",
INIT_33 => X"17400F7FBD75450800174AAFFD1555FFA2AA800105504001EFFFD140145557BE",
INIT_34 => X"0000000000000000000000000000000000000000000000020005D2E800BA0804",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000033FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"0405D434003F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"50805AC31007D6125724029216554A9847669903D640EC8E2001002604503004",
INIT_05 => X"07008000E0EA11803850C800010022660C1C0065003C0404002646DC20A02D40",
INIT_06 => X"30A03A0A138900001127A09234C81FF040000000002C44D620F0228454C83810",
INIT_07 => X"405584280B10014003A8067400920810FF3C72024300A0030048221ACEE383E4",
INIT_08 => X"1000C983E6041505253500F66E620428000B1804000152E52801A20200840900",
INIT_09 => X"0820500B90419005B0C309402030060860E01004A828408800440405E3502940",
INIT_0A => X"A2020010100007865421432121804021C20452880C2D200000045C18C0E0000A",
INIT_0B => X"371097006026226495446E2110AE4417411204400000306B8186185C42900693",
INIT_0C => X"A00308003080030800308003080030800308001840018400400602A018809800",
INIT_0D => X"4008081010108003C000210020460801001FB3650C50DB13111C0D95C20C2030",
INIT_0E => X"14804032007E281F840C00284A17210001060D8306C18360C1380A0260CB9808",
INIT_0F => X"1555D5D79BBEF8E50B041029075982BF3873041029079982BF39748AA0AC8000",
INIT_10 => X"5156AEA479BFD7F7F3041029075982BF3E73041029079982BF3F632C5F96D3C1",
INIT_11 => X"932C5F96A595405FC7F1CFEBC7586C4100A53162B47FD7E39FFEECE159870234",
INIT_12 => X"39464006FE037ACFB88083A99E06271BB0CA207DFDD5920057E0B001B0EBCC79",
INIT_13 => X"6F5DF5CA2A002DD51B6F7FC4A411D1E8D44517F14EAFE36E55150016EA8DB73E",
INIT_14 => X"9DB84953C30351452A13D55CFFA76E928E3891F148B30399F5FB7F28C800DFA0",
INIT_15 => X"110155AC57DFEAEF1005475F1D1F608819CF0EE76E12C824ADD9089715F25FAF",
INIT_16 => X"0D8360D834041A41A0000010180C02801680460FC900052FA10DC0006DA4881C",
INIT_17 => X"D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D836",
INIT_18 => X"8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360D8360",
INIT_19 => X"B000000000000000000000000020D8360D8360D8360D8360D8360D8360D8360D",
INIT_1A => X"1451451451448982C8A82E0820825942495377D9D701DC2E784601F8D187BEF8",
INIT_1B => X"4A2512A954AA5528944A25555145145145555555145145145555555145145145",
INIT_1C => X"FFC00000944A25128944A25128944A25128944A25128944A25128944A2512894",
INIT_1D => X"A5D2E820BA550000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFBFDFEFAAD142010007BEAB55FFAA821FFFFFFFFFFFFFFFFFFFFF7FBD74A",
INIT_1F => X"1FF002A821FFFFFFFFFEFF7D16AB55A2D542000A2D5400BA0800021FFFFFFFFF",
INIT_20 => X"DFFFFFFFC0010F7842AA10F780021FFFFFBFDF45A2D56AB45FFFFD54BAFF8000",
INIT_21 => X"6AB45A28000010082A975EFA2D140145007BC21FF5D2AAABFFF7D168B45AAD57",
INIT_22 => X"BC214555003DE10A2FBEAA00000002010552E95410AAFBD75FF5D7FEAB550051",
INIT_23 => X"04174AA5D00020BA555542145A284155FF5D517FE000004020AA552E80000F7F",
INIT_24 => X"00000000000017400082E954AA0800154AA0855575FFAAD57FE005D7BD740008",
INIT_25 => X"FFFFFDFEFF7FFD74AA552A820AA490A000000000000000000000000000000000",
INIT_26 => X"A080A051FFFFFFFFFEFF7F1FAFD7A2D5400001C7BEDB7DEBA4871FFFFFFFFFFF",
INIT_27 => X"6DFFFBD54AAE38E021FF0824821FFF7F1F8FC7EBD568B7DB6DF47000AADF400A",
INIT_28 => X"BC7E3D56AB7DB6DF78FD7EBF1C2000F78A2DA38E38A021C7E3F1F8F55AADB6FB",
INIT_29 => X"25EF497FEAB7D145B6FB45AA8E070281C20925FFBEDB451451C7BC01EF4124AD",
INIT_2A => X"00092412A87010E3F5C0145410E3DE28B6FFE8A101C0E05010412495428AAF1D",
INIT_2B => X"B7AE385D7FD74381400124825D0A000BA555F47145BE8A105EF555178E381C0A",
INIT_2C => X"00000000000000000000000000000154280024924AA1404174AA0055505EFBED",
INIT_2D => X"A80155FFFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA082A8000000000000000",
INIT_2E => X"F7FBD5410AAFBC00AA002A955FFF7FBFDFEFFFD568B45AAD5400005D7BFFFEFA",
INIT_2F => X"5AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF0000021EFF7D16AB55A2D56ABEF",
INIT_30 => X"45557BC21FF08003FF55AAD168BFFF7FFEAB45AAD140010F7AABFEBAAAAA8214",
INIT_31 => X"4100000154AAA2D1421FF007BE8BFF557BFDF55A2AA974AA5D04001EFFFFFD55",
INIT_32 => X"01EF55516AAAA5D2A82000082E95400A2D542155002ABDEBAF7FBE8A00552E95",
INIT_33 => X"174AA0855421FFFFFBEAAAA5D7BD74BA5D0002010552E820AA5D7BD7545F7AA8",
INIT_34 => X"0000000000000000000000000000000000000000000000174BA0004000AA5500",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000001000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000008128000000000000000000000024001620280000000000354200004008",
INIT_04 => X"000058800004C4024024001210001054B1C822009640000E2000002604003000",
INIT_05 => X"07008000E0200000000000000000200604000000001C04000026400000002C40",
INIT_06 => X"000000000000000004C010B35420015040000000002C42010010200004C83810",
INIT_07 => X"06E200201C00A14080082B26208008A009001201014022404402800408408020",
INIT_08 => X"00004180261C81210031000004340000200008105428020568040213003499C0",
INIT_09 => X"0000000990000000B0C308000000000860200160000000000038380000000000",
INIT_0A => X"10000000000005860000000080A0002060204080000000000004540800000000",
INIT_0B => X"00000000000000020001000022000000000000000000178000F8000101259000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000108000EC000000000000000010004B200000000000000000000000000",
INIT_0E => X"2000000000062801800400000000000000000000000000000000000000000000",
INIT_0F => X"828008084451B81A70AB3006BA0011400760AB3006BA0011400680F020968348",
INIT_10 => X"30B8011204082248A0AB3006BA0011400160AB3006BA0011400084C780687DBA",
INIT_11 => X"64C78068796E80A00802301BC0A7531EDD98E73B02800804620D030F873EB49F",
INIT_12 => X"B0A936B00000002044F091A860700FF9198AA115D5DA37F7A80C8A3604001C06",
INIT_13 => X"0000098551AC9000000000314E01F9F30198600631448410A2A8D64800000081",
INIT_14 => X"1046B2E00303842281C80A23004411AD661891F15148A4420804241526D60000",
INIT_15 => X"66A4A9D335F3D282000C6C5456C84850F61050C411AD6284FDA861682805A04A",
INIT_16 => X"0000000000000000000000000000000000004600C00138000030880042023043",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"9000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0C30C30C30C3451046260A9A69A603924554117747E18E0218CC01400163A20C",
INIT_1B => X"26934984C26130984C26130C30C30C34D30C30C30C30C34D30C30C30C30C30C3",
INIT_1C => X"FFC000004C26130984C26130984C26130984C26130984C26130984C26130984C",
INIT_1D => X"A5D2A800105D2E80000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFF7FBD74AA5D2E820BA55003DFFFFFFFFFFFFFFFFFFFFFFFFFD54A",
INIT_1F => X"B55FFAABDFFFFFFFFFFFFFFFFFDFEFF7FFD54BA5D2EA8BFFFF84021FFFFFFFFF",
INIT_20 => X"8B55A2D540010007BEAABAA2AE821FFFFFFFFFFFFFFBFDFEFAAD142010007BEA",
INIT_21 => X"021FFFFFFFFFEFF7D16AB55A2D542000A2D5400BA08003DFFFFFFFFFFFFF7FBE",
INIT_22 => X"FD54BAFF80001FF002ABDFFFFFFFFDFEFA2D56AB45AAFBD74AAFFD5420100804",
INIT_23 => X"FBE8B45AAD568BFFF7FBD74BAFF802ABFFFFAE821FFFFFBFDF45A2D56AB45FFF",
INIT_24 => X"0000000000002ABFFF7D168B45AAD57DFFFFFFFC0010F7842AA10F780155FFF7",
INIT_25 => X"FFFFFFFFFFFFBD54AA5D2A80000412A800000000000000000000000000000000",
INIT_26 => X"7E384071FFFFFFFFFFFFFFFFDFEFF7FFD74AA552A820AA490A38FFFFFFFFFFFF",
INIT_27 => X"D7A2D5400001C7BEDB7DEBA4BAFFFFFFFFFFFFF7FBFDFD7EBF1D24AA5D2AADBD",
INIT_28 => X"FFFFFFBFDFC7E3F5EAB45AAD140000007FEFA92A2AA851FFFFFFFFFEFF7F1FAF",
INIT_29 => X"74AAE3DF400000004021FFF7F1F8FC7EBD568B7DB6DF47000AADF400AA080A3F",
INIT_2A => X"F8F55AADB6FB6DFFFBD54AAE38E021FF0824BDFEFE3F1F8FD7AAD16DB7DBEFBD",
INIT_2B => X"A2DA38E38A125C7E3F1EAB55B6DB6FBD7E3F5D04AAFF8A2DBD7E3A0821C7E3F1",
INIT_2C => X"000000000000000000000000000002DBC7E3D56AB7DB6DF78FD7EBF1C2000F78",
INIT_2D => X"82AA8BFFFFFFFFFFFFFFFFFFFFF7FBD54BA552A80010002A8000000000000000",
INIT_2E => X"A2D5400AA552ABDF55A280155FFFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA0",
INIT_2F => X"FF7FBFDFEFFFD568B45AAD5400005D7BFFFEFAA8028BFFFFFFFDFEFF7FFFFF55",
INIT_30 => X"10AAFBC00AA002ABDFEFF7FBFDF55AAD16AB55AAD140010007BFFE10AAAA955F",
INIT_31 => X"B45A2D57DFFFFFFFD54AAA2FBC20100800021EFF7D16AB55A2D56ABEFF7FBD54",
INIT_32 => X"FF45AA8002145AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF00003FFEFA2D56A",
INIT_33 => X"EAB45AAD140010F7AABFEBAAAAA82155AAD568B55FFFFFDF55A2D1400AAF7AAB",
INIT_34 => X"00000000000000000000000000000000000000000000003FF55AAD168BFFF7FF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000002000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"000079800014CC02C034001600000000000000101EC0012EE0C0026E1E80F000",
INIT_05 => X"1F0FF433EFF0440C3902100002203F2EFC040388137C3E20C8EEC00284033CC0",
INIT_06 => X"7000660016490201700000000002FF57C8E8840155FDC0000010E40087D8787A",
INIT_07 => X"4000040007700000000000000001080FF900160000000200C00080001840BFE4",
INIT_08 => X"0009FFBFE5181606000410A4000004202AA8043E0000000000000001209244C0",
INIT_09 => X"0001227FB0000000F7DF78020004011FEFE00000000020031502000083880200",
INIT_0A => X"00000000000015BE0000004000000100000100506002008C2007D5FC80000024",
INIT_0B => X"0020000000000000000000000000000000210018800000000000000010000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000020",
INIT_0D => X"0008000000100000010000002000080101FFB600000000000000000000000000",
INIT_0E => X"0000003007FE29FF800C00000001002040000000000000020480002E42429C00",
INIT_0F => X"000000004D4E180010040000400000001E60040000400000001E6010003C0000",
INIT_10 => X"04000000000094B1E0040000400000001E60040000400000001E608040000004",
INIT_11 => X"0080400002000000000033628000100100000004000000006170C00080010000",
INIT_12 => X"B0020000000000295810000000A100020614148002000000000004307CC3CC00",
INIT_13 => X"000525802000000000014AC000120200000000003F0D800020100000000000A4",
INIT_14 => X"000020020C0C00000000002E2D000001006204040000000005786C0040000000",
INIT_15 => X"004000100A0C0939BEE1810080200000E0CE0EC000010020000000000000AE8A",
INIT_16 => X"000002008040400400C08080000000000049F6FFC01000000000000080080080",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"6902001000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"186186186190324C1090D0F3CF3CD039A060000600704000201120AB02090082",
INIT_1B => X"0C86432190C86432190C86596596596596596596596596596596596596596186",
INIT_1C => X"FFC00002190C86432190C86432190C86432190C86432190C86432190C8643219",
INIT_1D => X"A552A82010080400000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD54AA5D2A800105D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"0BA5500001FFFFFFFFFFFFFFFFFFFFFFFBD54BA552A8001000003DFFFFFFFFFF",
INIT_20 => X"FFEFF7FFD74BA552E801FF002E821FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E82",
INIT_21 => X"BDFFFFFFFFFFFFFFFFFDFEFF7FFD54BA5D2EA8BFFFF843FFFFFFFFFFFFFFFFFF",
INIT_22 => X"142010007BEAB55FFAA801FFFFFFFFFFFFFFBFDFEFFFD542000082EAAB55AAAA",
INIT_23 => X"FFFFFFFF7FBFDF55AAD140000087BE8B55F784021FFFFFFFFFFFFFFBFDFEFAAD",
INIT_24 => X"0000000000003DFFFFFFFFFFFFF7FBE8B55A2D540010007BEAABAA2AE975FFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA552A820001400000000000000000000000000000000000",
INIT_26 => X"81C0038FFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2A80000412ABFFFFFFFFFFFFF",
INIT_27 => X"EFF7FFD74AA552A820AA490A021FFFFFFFFFFFFFFFFFFEFF7FBD74BA5D2A8002",
INIT_28 => X"FFFFFFFFFFFFFFFBFDFEFFFFFD54BA5D2A801C7142E871FFFFFFFFFFFFFFFFDF",
INIT_29 => X"0010142AAFB7DBEAEBAFFFFFFFFFFFFF7FBFDFD7EBF1D24AA5D2AADBD7E38438",
INIT_2A => X"FFFEFF7F1FAFD7A2D5400001C7BEDB7DEBA4871FFFFFFFFFEFF7FBF8FD7E3D14",
INIT_2B => X"FEFA92A2AA925FFFFFFFDFEFE3F1FAF45A2D142010087FEDB55F78A051FFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFBFDFC7E3F5EAB45AAD140000007",
INIT_2D => X"02ABFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005D040000000000000000",
INIT_2E => X"F7FFD74AA5D2A800BA550428BFFFFFFFFFFFFFFFFFFFFF7FBD54BA552A800100",
INIT_2F => X"FFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA082A821FFFFFFFFFFFFFFBFDFEF",
INIT_30 => X"AA552ABDF55A2802ABFFFFFFFFFEFF7FBFFFFFF7FBD74BA552A80145552E955F",
INIT_31 => X"FEFF7FFEAB45AAD1420105D2ABFFFFFFAEA8BFFFFFFFDFEFF7FFFFF55A2D5400",
INIT_32 => X"DF55F7AE955FFF7FBFDFEFFFD568B45AAD5400005D7BFFFEFAA80175FFFFFBFD",
INIT_33 => X"6AB55AAD140010007BFFE10AAAA821EFF7FBFDFFFAAD168B55A2D542010007BF",
INIT_34 => X"00000000000000000000000000000000000000000000003DFEFF7FBFDF55AAD1",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"084A76341244919000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"000079800014CC03C075161E001118653D2408041FC004AEF000816E1C11F541",
INIT_05 => X"3F0F807BFFE000240100004683103E7FFE02482553FC3C0204EFC25010143CC0",
INIT_06 => X"1100441004201014B1709C910102FF5FC0A0000101FFE4036450E08247F87870",
INIT_07 => X"08750504800680102542AD800504530FF9061E8026998E9A00402CC25BD0FFFC",
INIT_08 => X"0011FBFFE04691A5A00101818A6800088228000001A044C8168480D010F200AA",
INIT_09 => X"B6E85A7FF080AC70FFDF78220010841EFFE7116E144071268DFD3E4C24040100",
INIT_0A => X"3151518A8A31B7FE00040009814C089202225412115428C03BC7D7FC15025B1A",
INIT_0B => X"1B1883007104032901CC63410ABD249C4B338934404037FC8BFE18008083B444",
INIT_0C => X"D9228D9228D9228D9228D9228D9228D9228D99146C9146C84006309044081A00",
INIT_0D => X"48000201800500941044312000900D4621FFBE00080081529904595123203040",
INIT_0E => X"308162029FFEADFF8050250010030165290008800440022201082401A002000C",
INIT_0F => X"5001318048A004A6C0D2820302C005A83480D1820302A009B02B101390C0CB28",
INIT_10 => X"485101408904831400D1820302C005A83480D2820302A009B02B021A85C09411",
INIT_11 => X"FA1A85C08834600024D052C1051E0B92D400360520202682C19024B6164E3004",
INIT_12 => X"C1B0D6404093E22A2012418A9D1D44ADD9E0F174103820101C0B8160D5516259",
INIT_13 => X"6C88660D8AA288209E615100280DA0052000C5006402000206C55144104D510C",
INIT_14 => X"024500A0D50020C04023033C52009144231D902818100C90058010361AC80812",
INIT_15 => X"198A12202386454988140600C0181500A13E830011008B0374007000B4E0CD00",
INIT_16 => X"008020080224004002000000703804008001F7FFF01B982B01258088C008CC41",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200802",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"F000000000000000000000000020080200802008020080200802008020080200",
INIT_1A => X"7DF7DF7DF7DFFFFEFEFFFE79E79FFFF3BC1FF3FDDFEFFFBEFFE7DF84081EFEFB",
INIT_1B => X"FEFF7FBFDFEFF7FBFDFEFF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF",
INIT_1C => X"FFC00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_1D => X"A5D2E80010000400000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA552A8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"0105D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E80010552EBFFFFFFFFFFF",
INIT_20 => X"FFFFFFFBD54BA5D2E82010002ABDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A80",
INIT_21 => X"001FFFFFFFFFFFFFFFFFFFFFFFBD54BA552A800100000001FFFFFFFFFFFFFFFF",
INIT_22 => X"BD74AA5D2E820BA5500001FFFFFFFFFFFFFFFFFFFFF7FBD74BA5D2E800BA5D00",
INIT_23 => X"FFFFFFFFFFFFFFEFF7FBD74AA552A800BA5D2E821FFFFFFFFFFFFFFFFFFFFF7F",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFEFF7FFD74BA552E801FF002E975FFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E800000800000000000000000000000000000000000",
INIT_26 => X"05D2ABFFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8200014003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFBD54AA5D2A80000412ABDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2E8000",
INIT_28 => X"1FFFFFFFFFFFFFFFFFFFFF7FBD54BA552E82028002AB8FFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74AA5D2E800AA5500021FFFFFFFFFFFFFFFFFFEFF7FBD74BA5D2A800281C0000",
INIT_2A => X"FFFFFFFFFFDFEFF7FFD74AA552A820AA490A071FFFFFFFFFFFFFFFFFFEFF7FBD",
INIT_2B => X"A801C7142E955FFFFFFFFFFFFFFFFDFEFF7FFD54BA5D2E80082492E871FFFFFF",
INIT_2C => X"0000000000000000000000000000038FFFFFFFFFFFFFFFBFDFEFFFFFD54BA5D2",
INIT_2D => X"D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008000000000000000000",
INIT_2E => X"FFFBD54AA5D2E800005D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFF7FBD54BA552A80010002ABDFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"AA5D2A800BA5504021FFFFFFFFFFFFFFFFDFEFF7FBD74AA552E820BA002AA8BF",
INIT_31 => X"FFFFFFBFDFEFFFFFD54BA552E800BA5D04021FFFFFFFFFFFFFFBFDFEFF7FFD74",
INIT_32 => X"0000082A955FFFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA082A955FFFFFFFF",
INIT_33 => X"FFFFFF7FBD74BA552A80145552E975FFFFFFFFFEFF7FBFDFFFFFFBD74AA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000002ABFFFFFFFFFEFF7FB",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"431965109E4481D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"492C0020220001010E4916C884DCD607E5EC2A344103E48003D0800023D0072C",
INIT_05 => X"00107C441001100D620A06D683018001023D37E5088043620101179092540112",
INIT_06 => X"401002010042384D223C19C3552800081ADA0E054402365774611E047020008E",
INIT_07 => X"491EC04ED017AB5497EB923F08182E20020689B735011FBFE7BC062602944019",
INIT_08 => X"154A00401D4425ADA9035BE19C8F9442A8801200F4C9D7AC8093A051727B2AC3",
INIT_09 => X"9A50020040E48D50080002B00A0C00801014541E9504703680017F6CB4050700",
INIT_0A => X"8151538A8A738041C23020131A80CFDFF3FE509A907C6AC05040220409009031",
INIT_0B => X"2D040050110081E9528963546278008AA80381B4000500026800000109379864",
INIT_0C => X"1C2A81C2A81C2A81C2A81C2A81C2A81C2A81C9540E1540E00140000610000320",
INIT_0D => X"594A06870A9CA0D458D131652A154D46B6000850800801628013456520CA0928",
INIT_0E => X"02080448C00044000A1EC1C44140D101A54280A14050A028500A84F02842A24C",
INIT_0F => X"0061338359E0C4E6C256690581800F1C3E82562B0581200F1C3F081456022804",
INIT_10 => X"2C438100AB8581B602562B0581800F1C3E8256690581200F1C3F1238473F1210",
INIT_11 => X"2238473F0E1050083750B3E4275F829547008600C030374361FA2CEE046D4812",
INIT_12 => X"C1128C4CC012A66F61154C019511628756231018500C00203E13806156516078",
INIT_13 => X"54CDE608AA612C0096C37B00D1724801A0009C606D1221D104553096004B61BC",
INIT_14 => X"870B012A41E0F0600035842E7601C2C4AC68A98810080AA825A8902251899802",
INIT_15 => X"58234A89637E00D0A1080301401C390320188321C2C0B13890105800D520AF94",
INIT_16 => X"8822088222F110111B281A54753AA004002601001918008C10912A4440B24E8B",
INIT_17 => X"8220882208822088220882208822088220882208822088220882208822088220",
INIT_18 => X"2008020080200802008020080200802008020080200802008022088220882208",
INIT_19 => X"E82891448000000001FFFFFFFFC8020080200802008020080200802008020080",
INIT_1A => X"3CF3CF3CF3DFFBFEFEBEEEFBEFBEFBEBFDF7F7FBDFD1FE3EFBD7ADFBF7EFBEFB",
INIT_1B => X"FE7F3F9FCFE7F3F9FCFE7F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"FFC00001FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"A5D2E82000000000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8000008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74AA552E8000055003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A82",
INIT_21 => X"BFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E80010552EBFFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD54AA5D2A800105D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A82000552A",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD54AA5D2A800005D2EBDFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"000000000000001FFFFFFFFFFFFFFFFFFFFFFFBD54BA5D2E82010002AA8BFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100004000000000000000000000000000000000",
INIT_26 => X"008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA552A8200014003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E800105D043FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"54AA5D2A82010552EBDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2E800005D2ABF",
INIT_2A => X"FFFFFFFFFFFFFFFFFBD54AA5D2A80000412AB8FFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E82028002AA8BFFFFFFFFFFFFFFFFFFFFFFFBD54BA552E80038492EB8FFFFFFF",
INIT_2C => X"00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFF7FBD54BA552",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000040000000000000000",
INIT_2E => X"FFFFD74BA552A8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E800000",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005D043FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"AA5D2E800005D2EBDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA552E8001055003FFF",
INIT_31 => X"FFFFFFFFFFFFF7FBD54BA5D2A820105D2ABDFFFFFFFFFFFFFFFFFFFFFFFFBD54",
INIT_32 => X"00AA082EA8BFFFFFFFFFFFFFFFFFFFFF7FBD54BA552A80010002AA8BFFFFFFFF",
INIT_33 => X"FDFEFF7FBD74AA552E820BA002AAABFFFFFFFFFFFFFFFFFFEFF7FBD74BA552E8",
INIT_34 => X"0000000000000000000000000000000000000000000000021FFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"2C4360101A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"00017B810015DC03D034201E14000036486008101FC0002EE006297E1C05F561",
INIT_05 => X"BF0F817FFFE80100004044800080BEFFFC0248005FFC3C18A5FFC2444484BCC0",
INIT_06 => X"B0801408110000109127E0500002FFDFC000000001FFC0832050E00047F97870",
INIT_07 => X"00D1D72040048D00388387D03D0E591FFD201F862691DFBE077C2BC45B40FFE4",
INIT_08 => X"001FFBFFEC440501A5604B31062356282AA84200D12342113EDC400000045828",
INIT_09 => X"25A890FFF0002023FFDF79000000000EFFE309606020008005FC000000402000",
INIT_0A => X"30000000000037FF50010103134CAFDF03BA18000F39A0106F87D7FA84024B02",
INIT_0B => X"1B188300624483890564084198AD249C43300C00415037FC83FE1840C0902400",
INIT_0C => X"C1010C1010C1010C1010C1010C1010C1010C10086080860840063090442A1800",
INIT_0D => X"0001403000100200180480000095280001FFBF040C40C81119A41C1443243050",
INIT_0E => X"32A163821FFEAFFF805025E00853B92588000400020001000020A80180080020",
INIT_0F => X"90401486148484054395E27E428002A4200397E07E422002A420100382FCC308",
INIT_10 => X"641100C0788417000397E07E428002A4200395E27E422002A420110A51C01C05",
INIT_11 => X"C90A51C01A2490040590C08120558C1759BE1C05A0400383808800DA1929F728",
INIT_12 => X"00CE720000136006000215EA0A4833A32C8832050028603050014031B3950000",
INIT_13 => X"6C00C006658280009A2030108B14AC05C00112405222088B8332C140004D1018",
INIT_14 => X"A2659196B6808060201281004228996085F10020180C030880D11019CE400002",
INIT_15 => X"0108152A49DC7143F01C04240030720641E0A028996483A17204680410A04104",
INIT_16 => X"040100401000080080000000000002001201F7FFC0011C2F81A48080CA32800A",
INIT_17 => X"4010040100401004010040100401004010040100401004010040100401004010",
INIT_18 => X"0100401004010040100401004010040100401004010040100401004010040100",
INIT_19 => X"0000000000000000000000000000401004010040100401004010040100401004",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000020000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFC0000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2A8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E80",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8000008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA552A8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A820000004",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA552A8201000043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E8000055003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA552A8200008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001008043F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA552A8200014003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E800105D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E820101C003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552",
INIT_2D => X"0043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA552A8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001008043FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74AA552A8200008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"200055043FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005D043FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD54AA552E8001055003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA552E8",
INIT_34 => X"00000000000000000000000000000000000000000000003DFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"00003A2E200811000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"000079800014CC03C034001E04010850300000101FC0002EE000006E1C00F500",
INIT_05 => X"1F0F8033FFE000000000000000003E2FFC024800137C3C0000EFC00000003CC0",
INIT_06 => X"000000000000000091C115500002FF5FC000000001FFC0000010E00007F87870",
INIT_07 => X"10E600084002040A10812A000500590FF9001F95406A8000037230C01840FFE0",
INIT_08 => X"0001FBFFEC4695A501604A000C7585080002C200408102F16C0184800026C92C",
INIT_09 => X"24A8107FF0000000FFDF78000000000EFFE001600000000005FC000000000000",
INIT_0A => X"30000000000037FF4000000AA0354000019C4000012800002387D7F804024B02",
INIT_0B => X"1218830060040A04000400000801241443300800404037E883FE180000000000",
INIT_0C => X"C1000C1000C1000C1000C1000C1000C1000C1000608006084006301044081800",
INIT_0D => X"00000004800B0000000000000000000001FFBE00080080101904181003003000",
INIT_0E => X"B08062021FFEADFF800020800000002088000000000000000000200180000000",
INIT_0F => X"D0210840009181008024A00043601100210024A00043C0110020901382CCCB28",
INIT_10 => X"0C920180040A03080024A00043601100210024A00043C01100209240C840C201",
INIT_11 => X"1A40C840A604E0080820009908008341B000A821207008200289001006832086",
INIT_12 => X"0166B40600800082041205EC00044C1ACB66C37542082030281E058000101281",
INIT_13 => X"0010480B27A004300004103160DB3005E000618040C022000593D00218000209",
INIT_14 => X"880012BBFF20406040084210C062000C2A2DDD00180C04504086002CD680C010",
INIT_15 => X"4106020804295C98F80400008040CC0582169022000C2876C404780028500160",
INIT_16 => X"000000000000000000000000000000000001F7FFC001B823018F008800088052",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"C800000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"7CF7CF7CF7D933CC3090CABAEBAFF969319815DD5EDCF9822659AE7B095A220C",
INIT_1B => X"1E0F0783C1E0F0783C1E0F7DF7DF7DF3CF3CF3CF3CF3CF7DF7DF7DF7DF7DF7CF",
INIT_1C => X"FFC000003C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C",
INIT_1D => X"A5D2E82010080400000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"00000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E800000800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8001000003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100804000000000000000000000000000000000",
INIT_26 => X"000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"A8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000043FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008040000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8000008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"000008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2A8001008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00002000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"924279824C94CC1BE0B4001F20000000020380401FE0082EF000106E1C00F500",
INIT_05 => X"1F0F8033FFF048202582800100523E2FFE024820137C3C0040EFE02000003CE4",
INIT_06 => X"F10466105670019C900000100002FF5FC0E0801101FFC0000010E08A07FC7870",
INIT_07 => X"0000040000000000000000000500590FF9001F0000000000033020C01840FFFC",
INIT_08 => X"0001FBFFFD0004000100502000011400000282004001020000000001009015C0",
INIT_09 => X"2CB8DA7FF8004000FFDF7C062031863EFFF75D78004001010DFC000020050100",
INIT_0A => X"30000000000037FFC00602000000000001980400002800032387D7FE94FBEF2B",
INIT_0B => X"9258830060040200000400000801243443B00808404037E883FE180C00000000",
INIT_0C => X"C1000C1000C1000C1000C1000C1000C1000C10006080060840077330C4889CC2",
INIT_0D => X"0000000000000000000000000001280001FFBE00080080101904189003003000",
INIT_0E => X"30A063021FFEADFF805025C0304001E58906088304418222C108A009A0904000",
INIT_0F => X"1000000000100100000480000200100000000480000200100000100380F0C308",
INIT_10 => X"0010000000080000000480000200100000000480000200100000000040400000",
INIT_11 => X"0000404000040000000000080800000110000000200000000200000000012000",
INIT_12 => X"00021000000000800002018C0100000208000008001220000000040040000080",
INIT_13 => X"0010000020800000000400000010200200000000008002000010400000000200",
INIT_14 => X"0800000210000080010000008002000000210000201000000002000042000000",
INIT_15 => X"0184000000084000000006050000000002000002000000204000000000000020",
INIT_16 => X"08822288226410410346010000000400A011F7FFE00318230104008000008000",
INIT_17 => X"8822088220882208822088220882208822088220882208822088220882208822",
INIT_18 => X"8220882208822088220882208822088220882208822088220882208822088220",
INIT_19 => X"0404000017FFFFFFFFFFFFFFFFE0882208822088220882208822088220882208",
INIT_1A => X"492082492085048029890AD34D35FDD04A165129432D518B45265EFC30760AED",
INIT_1B => X"C46231188C46231188C462492492492492492492492492082082082082082082",
INIT_1C => X"FFC000058AC562B158AC562B158AC562B158AC562B158AC562B158AC562B158A",
INIT_1D => X"A5D2E820100800000000000000000000000000000000000000000000000003FF",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100000",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000043FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"4A53D958C50000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"DBFAFBD7FB1CDEBEF1BE17F7AC88042787FBFFF8FEE9FF7EE6F4C0EE1FFAF869",
INIT_05 => X"5F0FFEB3EFFEFFBDA7F7FED508707E2EFEBF6FFEB37C3FF302EEEDFF9B487CF6",
INIT_06 => X"74EADE4EBDFDAC9930F6F8129E3FFFF7C3E3A74667FDDB7FB870FF30FFDEF87F",
INIT_07 => X"8173840C07783060C72DF7D828912E6FFB80162776F3BFB7077E82255E40BFEF",
INIT_08 => X"4769FFBFE43C872321367036163F1C0820A3063F460D1AEFC000060042648C41",
INIT_09 => X"BEFB967FBD13D981F7DF7D7E6171AF3FEFE8A3E679FAC1FD1FFFBEB000763A84",
INIT_0A => X"F3A3AD1D1DAD7FBE7D67D7F3BB79CFFB83BF14EC1E7D7300B017F5FFE6FBEF73",
INIT_0B => X"52199F58F6EE6F5E7FAC4C03DB856CD4CF720FE8C4427FF8CFFE38FF7F6BD928",
INIT_0C => X"F78C0D78C0D78C0D78C0D78C0D78C0D78C0D7A606BC606B8C56F7730ECCDBDF1",
INIT_0D => X"EA035CF6100C0E60FB9FC3A80EF69A04DFFFF7FF5E75FF341B867D3683A03A40",
INIT_0E => X"36B867027FFFF9FF8FAFAA3ADEBFB9726BAF5FD7AFEBD7F7EFFD7ACDB7F947F0",
INIT_0F => X"10003E020080A40403E8BD8002000FC02003E8BD8002000FC02010979AFFE36C",
INIT_10 => X"80100000EE00034003E8BD8002000FC02003E8BD8002000FC020037B0040A000",
INIT_11 => X"037B0040C00400003D80008160400FD81341C00020003B80008C00801EF02853",
INIT_12 => X"01F1190981038406809677FA080468C46A81080581002000780C8001C8100201",
INIT_13 => X"7080D00F90D162001C803411FC0024080001F80040026C0807C868B1000E401A",
INIT_14 => X"B02013F810503A00003E020042AC080CEB01228A80000F600080123E23213040",
INIT_15 => X"61F810087520750001064180807868000110C02C080CFA0042400000F8800105",
INIT_16 => X"5FD7F7FDFF7EFEEFF3EEC3FF7FBFFBCB7FFFFEFFE00BFF7FEBF420800EC0CBEE",
INIT_17 => X"FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F",
INIT_18 => X"D7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5",
INIT_19 => X"6DAE443237FFFFFFFFFFFFFFFFF5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5FD7F5F",
INIT_1A => X"4D34D30C30DD795EAA6AFC38E38EA3AB788962B79E923C2CD990A7D3B4A9FC37",
INIT_1B => X"26130984C26130984C26130C30C30C30C30C30C30C30C30C30C30C30C30C30C3",
INIT_1C => X"FFC000004C26130984C26130984C26130984C26130984C26130984C26130984C",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"0842D85841000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"DBEAE5D6D91C2EBCE1B21EA72C00000007FBE7C8F8E9EF79E6D440E91FDAE061",
INIT_05 => X"5C8FFCB38FF6B68984B5BCE408347E28FEBF6FEEB3723F7102E8EDBF8A4872F6",
INIT_06 => X"946ACF46ACE0841A00006A089E3FFF27C3032646EFF1DB7FA868FE30EF1CE47E",
INIT_07 => X"8000000A20083060C00C81882A008C6FF880060424B39FB6037F00051C003FE0",
INIT_08 => X"4761FA3FE4010440410844060001040A00002200460D1A060000050400000010",
INIT_09 => X"FEEB027E390A4881C7BEFC5F6171CE2F8FE823E778DAC16C1FFBBC9000315895",
INIT_0A => X"F606013030213C3E2D62D6E21259CFDB039E806C024531008017C1F826FFEF41",
INIT_0B => X"5219AB5AF86F7D5E382A440349816DD4C7560B60D4427FF0C7FEBABF3F6BD108",
INIT_0C => X"E3440C3440C3440C3440C3440C3440C3440C3C2061A2061AD46FF730E5CCBCD5",
INIT_0D => X"6203E8FC10080A20ED1D41880CC61A044DFFC6EB5AB5B7941BC63F1683803C00",
INIT_0E => X"B88572023FFE91FF98AEAA1AC6AC9A3A4AAD5B56ADAB56D5AFD572C597B14750",
INIT_0F => X"10003E020000260403C8948002000EC0000BC8948002000EC00010878AC3CB8A",
INIT_10 => X"80100000EE0000400BC8948002000EC0000BC8948002000EC000097B00402000",
INIT_11 => X"017B0040400400003D80000070400DD81041400020003B80000410801AF02041",
INIT_12 => X"05D11101010384008086378A080428C46A80080081002000780C800188000301",
INIT_13 => X"7080102E909042001C800409FC0020080001F80000007C0807484821000E4002",
INIT_14 => X"F02003F810100A00003E020000BC0808EB01020280000F60000002BA22202040",
INIT_15 => X"21F810007520750000024080807868000100403C0808FA0040400000F8800001",
INIT_16 => X"5B56D5B5EF3AF6AF6389C2FE128971AB2DDDF8FFE0031B776BF4208006C0C926",
INIT_17 => X"B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D",
INIT_18 => X"56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B56D5",
INIT_19 => X"238B443A3FFFFFFFFFFFFFFFFFD5B56D5B56D5B56D5B56D5B56D5B56D5B56D5B",
INIT_1A => X"00000000000F0080397908000000A4805F09C42D0200903950C086D420010825",
INIT_1B => X"8040201008040201008040000000000000000000000000000000000000000410",
INIT_1C => X"FFC00005028140A05028140A05028140A05028140A05028140A05028140A0502",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100804",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"461080404900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"00800040110102000902002000888400081045A8A00003C00000500000080008",
INIT_05 => X"0000000000024CA0A0101800032000400000000B800000014000000B08180000",
INIT_06 => X"0020280202802C00020800008A14002011110012220009A88800009A88000000",
INIT_07 => X"8108044200091224484510201000204000800020410000000080000104000009",
INIT_08 => X"132800000140200808021006108010422AAA8000224489028492201140092240",
INIT_09 => X"0001C800004080A0000002480B04008100011000088800081002C19020150B00",
INIT_0A => X"4353529A9A528000040040702080000000400064080011001050000200000018",
INIT_0B => X"01400048012220122A0004168110400004000040811600000400001036584108",
INIT_0C => X"36050160501605016050160501605016050160280B0280B00120008430660210",
INIT_0D => X"2A000C4210040860B188C0A8065302005A0040390010120500002002C0040010",
INIT_0E => X"8221050060001000028000080205001066000100008000400490020402010530",
INIT_0F => X"000000000000A00000081480000001400000081480000001400000800C010820",
INIT_10 => X"8000000000000240000814800000014000000814800000014000000100002000",
INIT_11 => X"000100004000000000000001400000080041400000000000000C000000100041",
INIT_12 => X"000101010100000480802A400000004000000800810000000000000048000000",
INIT_13 => X"0000900010104200000024000400000800000000000244000008082100000012",
INIT_14 => X"1000004000100A00000000000284000040000202800000000000120020202040",
INIT_15 => X"2050000010000000000240800000000000104004000040000040000000000005",
INIT_16 => X"010040108408420430E699AA42A1508104EA08000000810020000000044001AC",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"0506117080000000000000000000100401004010040100401004010040100401",
INIT_1A => X"4104104104006C1A8283AC618618EF10C0422205822140048D2E581E80DEC4D2",
INIT_1B => X"C06030180C06030180C060410410410410410410410410410410410410410410",
INIT_1C => X"FFC0000582C160B0582C160B0582C160B0582C160B0582C160B0582C160B0582",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"00000003FFFFFFFFC00000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0401D940CD0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"49B87A417315D20A313E17F1800000058013DDF8BE21F36E02F0D06E03E8F800",
INIT_05 => X"1F007E33E01A4D9C87525E5101603E6E023D27DA937C03E340EE25CB9B483C12",
INIT_06 => X"F0A05A0A15AD0C0130F6F0128A16FFF001E1870223FC3BFC98101F109FC6780F",
INIT_07 => X"8073800407781020476467D008910A4FFB80100332D1AE93059282215E408006",
INIT_08 => X"0221FF80003C832320342036063F08000001063F42050AEB4000221000248C01",
INIT_09 => X"9A51547F8C1111A0F041056A0100A11FE000916249A800B915FE82B020522900",
INIT_0A => X"42A2AD1515AD5780540541619968C76980E914E4163D53002017F405C409A42A",
INIT_0B => X"0140140816A22B126DA40C03531440800C2005C8800217F80C000055FF7C4928",
INIT_0C => X"268D0068D0068D0068D0068D0068D0068D006A68034680300021410028450530",
INIT_0D => X"AA01587410080C60AB0F42A804628200DBFFF13D04505B2500806522C0A40A50",
INIT_0E => X"941922006FFFF8000F8F80281A16A1504302058102C0816244B82A0CA25907D0",
INIT_0F => X"000000000080A40000283D80000001402000283D80000001402010901A7D6944",
INIT_10 => X"800000000000034000283D80000001402000283D80000001402002010000A000",
INIT_11 => X"02010000C000000000000081600002080341C00000000000008C000004100853",
INIT_12 => X"0021090981000006809076B20000404000010805810000000000000048100200",
INIT_13 => X"0000D0011051620000003410040004080000000040026C00008828B10000001A",
INIT_14 => X"B000104000503A000000000042AC00044000228A800000000080120421213040",
INIT_15 => X"607800081000000001064180000000000010C02C000440000240000000000105",
INIT_16 => X"05816258964C4A44A0C689FF3F9FFEC5D6DBFE0020096528A0B000000CC043EC",
INIT_17 => X"5816058160581605816058160581605816058160581605816058160581605816",
INIT_18 => X"8160581605816058160581605816058160581605816058160581605816058160",
INIT_19 => X"F506003017FFFFFFFFFFFFFFFFE0581605816058160581605816058160581605",
INIT_1A => X"5D75D75D75DFFFFEFCFDF7FFFFFF5DE7FC3DF3F2DDCFFFBEFFCF1F84421FFEFF",
INIT_1B => X"EFF7FBFDFEFF7FBFDFEFF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF7DF75D7",
INIT_1C => X"FFC00007DFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDF",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"E800000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"3CF3CF3CF3DD7FDEBAFAFEFBEFBFFBFBB9DFF7FFDFF3FC3EFFF7FDFBBDFFFEFF",
INIT_1B => X"FE7F3F9FCFE7F3F9FCFE7F3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF3CF",
INIT_1C => X"FFC00001FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"08425818000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"DB6A618248140C18E0B016872400000007EBA24058E1ECA8E2D400681FD0E061",
INIT_05 => X"1C0FFC338FF01009048084C400103E28FE3F6FE513703F7000E8E5B4825030F6",
INIT_06 => X"100046000460001800006800142AFF07C202060445F1F2572060FE82671C607E",
INIT_07 => X"00000008800020408008818838000C2FF800060424B39FB6037E000418003FE0",
INIT_08 => X"0441FA3FE4000400010040000001040880000200440912040000040000000000",
INIT_09 => X"BEE8027E38004801C79E7C162231862E8FE00166704041240DF93D0000000000",
INIT_0A => X"B00000000000343E002202021259CFDB039E0008024520000047C1F804FBEF01",
INIT_0B => X"121883107044094C1028400548812494C3120920404437F0C3FE180D89279000",
INIT_0C => X"C1000C1000C1000C1000C1000C1000C1000C18006080060840477330C4889CC0",
INIT_0D => X"400340B400080200481501000884080405FF86400800811019861D1403803800",
INIT_0E => X"308062021FFE81FF880EA000400098200C04080204010200810020C180904240",
INIT_0F => X"10003E020000040403C0800002000E800003C0800002000E8000100780C2C308",
INIT_10 => X"00100000EE00000003C0800002000E800003C0800002000E8000017A00400000",
INIT_11 => X"017A0040000400003D80000020400DD01000000020003B80000000801AE02000",
INIT_12 => X"01D01000000384000006118A080428846A80000000002000780C800180000201",
INIT_13 => X"7080000E808000001C800001F80020000001F8000000280807404000000E4000",
INIT_14 => X"A02003B810000000003E020000280808AB01000000000F600000003A02000000",
INIT_15 => X"01A81000652075000000000080786800010000280808BA0040000000F8800000",
INIT_16 => X"08020080223010010308025410082404A015F0FFE003182701B420800280C802",
INIT_17 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_18 => X"0200802008020080200802008020080200802008020080200802008020080200",
INIT_19 => X"0008004017FFFFFFFFFFFFFFFFC0802008020080200802008020080200802008",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"FFC0000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"A5D2E82010080000000000000000000000000000000000000000000000000200",
INIT_1E => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_1F => X"01008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFF",
INIT_20 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_21 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_22 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_23 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_24 => X"0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_25 => X"FFFFFFFFFFFFFD74BA5D2E820100800000000000000000000000000000000000",
INIT_26 => X"008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_27 => X"FFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201",
INIT_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_29 => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_2A => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_2B => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_2C => X"000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_2D => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000000000",
INIT_2E => X"FFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_2F => X"FFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFF",
INIT_30 => X"BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFF",
INIT_31 => X"FFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74",
INIT_32 => X"201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFF",
INIT_33 => X"FFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8",
INIT_34 => X"00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


end;