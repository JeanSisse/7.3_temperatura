library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_master is
	port(clk             : in  std_logic;
        address_a       : in  std_logic_vector(31 downto 2);
        enable_a        : in  std_logic;
        wbe_a           : in  std_logic_vector(3 downto 0);
        data_write_a    : in  std_logic_vector(31 downto 0);
        data_read_a     : out std_logic_vector(31 downto 0);

        address_b       : in  std_logic_vector(31 downto 2);
        enable_b        : in  std_logic;
        wbe_b           : in  std_logic_vector(3 downto 0);
        data_write_b    : in  std_logic_vector(31 downto 0);
        data_read_b     : out std_logic_vector(31 downto 0));
end; --entity ram     

architecture ram_master of ram_master is
signal enable_a_lo       : std_logic;
signal wbe_a_lo          : std_logic_vector(3 downto 0);
signal data_write_a_lo   : std_logic_vector(31 downto 0);
signal data_read_a_lo    : std_logic_vector(31 downto 0);
signal enable_b_lo       : std_logic;
signal wbe_b_lo          : std_logic_vector(3 downto 0);
signal data_read_b_lo    : std_logic_vector(31 downto 0);
signal enable_a_hi       : std_logic;
signal wbe_a_hi          : std_logic_vector(3 downto 0);
signal data_read_a_hi   : std_logic_vector(31 downto 0);
signal enable_b_hi       : std_logic;
signal wbe_b_hi          : std_logic_vector(3 downto 0);
signal data_read_b_hi    : std_logic_vector(31 downto 0);
signal address_a_reg     : std_logic_vector(31 downto 2);
signal address_b_reg     : std_logic_vector(31 downto 2);
signal enable_a_lo_256       : std_logic;
signal wbe_a_lo_256          : std_logic_vector(3 downto 0);
signal data_write_a_lo_256   : std_logic_vector(31 downto 0);
signal data_read_a_lo_256    : std_logic_vector(31 downto 0);
signal enable_b_lo_256       : std_logic;
signal wbe_b_lo_256          : std_logic_vector(3 downto 0);
signal data_read_b_lo_256    : std_logic_vector(31 downto 0);
signal enable_a_hi_256       : std_logic;
signal wbe_a_hi_256          : std_logic_vector(3 downto 0);
signal data_read_a_hi_256   : std_logic_vector(31 downto 0);
signal enable_b_hi_256       : std_logic;
signal wbe_b_hi_256          : std_logic_vector(3 downto 0);
signal data_read_b_hi_256    : std_logic_vector(31 downto 0);
begin
process(clk)
begin
if rising_edge(clk) then
	address_a_reg <= address_a;
	address_b_reg <= address_b;
	end if;
end process;
data_read_a <= data_read_a_lo when (address_a_reg < x"0001000"&"00") else
data_read_a_hi when ((address_a_reg >= x"0001000"&"00") and (address_a_reg < x"0002000"&"00")) else 
data_read_a_lo_256 when ((address_a_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_a_hi_256 when ((address_a_reg >= x"0003000"&"00") and (address_a_reg < x"0004000"&"00"));
data_read_b <= data_read_b_lo when (address_b_reg < x"0001000"&"00") else
data_read_b_hi when ((address_b_reg >= x"0001000"&"00") and (address_b_reg < x"0002000"&"00")) else
data_read_b_lo_256 when ((address_b_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_b_hi_256 when ((address_b_reg >= x"0003000"&"00") and (address_b_reg< x"0004000"&"00"));
enable_a_lo <= enable_a when (address_a < x"0001000"&"00") else '0';
enable_b_lo <= enable_b when (address_b < x"0001000"&"00") else '0';
enable_a_hi <= enable_a when ((address_a >= x"0001000"&"00") and (address_a < x"0002000"&"00")) else '0';
enable_b_hi <= enable_b when ((address_b >= x"0001000"&"00") and (address_b < x"0002000"&"00")) else '0';
enable_a_lo_256 <= enable_a when ((address_a >= x"0002000"&"00") and (address_a < x"0003000"&"00")) else '0';
enable_b_lo_256 <= enable_b when ((address_b >= x"0002000"&"00") and (address_b < x"0003000"&"00")) else '0';
enable_a_hi_256 <= enable_a when ((address_a >= x"0003000"&"00") and (address_a < x"0004000"&"00")) else '0';
enable_b_hi_256 <= enable_b when ((address_b >= x"0003000"&"00") and (address_b < x"0004000"&"00")) else '0';
wbe_a_lo <= wbe_a when  enable_a_lo='1' else x"0";
wbe_a_hi <= wbe_a when  enable_a_hi='1' else x"0";
wbe_b_lo <= wbe_b when  enable_b_lo='1' else x"0";
wbe_b_hi <= wbe_b when  enable_b_hi='1' else x"0";
wbe_a_lo_256 <= wbe_a when  enable_a_lo_256='1' else x"0";
wbe_a_hi_256 <= wbe_a when  enable_a_hi_256='1' else x"0";
wbe_b_lo_256 <= wbe_b when  enable_b_lo_256='1' else x"0";
wbe_b_hi_256 <= wbe_b when  enable_b_hi_256='1' else x"0";



ram_bit_0_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"88280C4C7B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"00160090920C04800904848262220277E05152B280780D407428E723C01E1400",
INIT_05 => X"0006D46207801E400183C0707800E6000E008057641E00473C40680D32330C00",
INIT_06 => X"C165000225E2C11E2C12A0D0144AC27206582C166504816162002000B0FC21D5",
INIT_07 => X"5E6D233B964E7CD99DFB870E1DDDD889C5FBDC440129A0604442180238203F70",
INIT_08 => X"AD23C17544C581000657A0E8E83D86F0E4A7B2D88AAAFD7FE0E1833AC5920CFC",
INIT_09 => X"6D82082E2081B6C0027ADA398000008A504318404005B70663212C04A080B036",
INIT_0A => X"414568729139FA5610C00001A2502440888420247041E87681008CE9AFC80001",
INIT_0B => X"22B826E250B12346F1244812240912048941621804A150CA1CA45C254D4AF4AA",
INIT_0C => X"F80FA97FE0F0009E0FC40FA97FE0F0009E0FC048211E9C11C31F82E4A0008900",
INIT_0D => X"040FAB3FE0F0009E0FC40FAB3FE0F0009E0FCC42EFDFBF0AE03080E2AEB2E0F1",
INIT_0E => X"013879BA878FE807F65FBF12E0380231F0BD9E3FC08FEBD6F661C0E008C3CB5F",
INIT_0F => X"B248831ACBFC8BBDCAB779BC699F20180309A0F83BE2B87C7C42EFDFBF187806",
INIT_10 => X"4131B59003FFEC07F00003F01FB90BE9F01FC8B38C2098DAE007F323A0C83136",
INIT_11 => X"3080E29F1B2BE9F8A27E6E915C0E004C72BEC800FE7464290626D7003F994718",
INIT_12 => X"FC0C2352A0024B83F07F198BE9F8A0FFDA2A3C0202B8776A2FA7F023F7D06570",
INIT_13 => X"1448126105810941C5C068000CD4004C0905E52630BB1AE49C2BA7F98D6F846D",
INIT_14 => X"6074EA560F0416A24844B01302A26100C4801844069B0C88881A28C141118000",
INIT_15 => X"A781E2781EA781E2781C33C0613C0E21020800239450116ED443C041B47E9665",
INIT_16 => X"241140A056954AB0C280D0002020187007122C3E04E03383E2781EA781E2781E",
INIT_17 => X"20481204812048120481204812048120481204812048120481204812058112C1",
INIT_18 => X"0481204812048120481204812048120481204812048120481204812048120481",
INIT_19 => X"0000000000001204812048120481204812048120481204812048120481204812",
INIT_1A => X"C4109CAF9C4C83B8E38E2AE9C136AD8E9B562CF042E6281CF13043A85D400000",
INIT_1B => X"F0F87C3E08208208208208208208208208208208208208208208208208208220",
INIT_1C => X"1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1",
INIT_1D => X"000000000000000000000000000000000000C3007FFFFFFFFFFFA00000F87C3E",
INIT_1E => X"4214555517DEAA5D7BFFEAAF7803FEBAF7FFD74BAAAAABDEBAF7AE8000000000",
INIT_1F => X"1555FF55517FE000055421FF00557DF45A2D5401EFF7D142145A2AE800BA0851",
INIT_20 => X"5555555A2AABFFFF5D516AA00A28028A00AAAEBFE00A2FBD75FFFF8400155085",
INIT_21 => X"5517FF45A2AEBDEBAAAAAA8BFFF7D140010FF84174BA552EBDFFF0004020005D",
INIT_22 => X"5504000BA5D2E97545A28028B4508554014508043FEBA082ABFE10AAAEA8ABA5",
INIT_23 => X"FA2AABFE00FFFFD74AA085540000002E801FF557FD75FF0051401FF5D0015410",
INIT_24 => X"EFF7FFC20BAF7D1575450800020BA08517FF45F7FBFFF45A2FFFDE00002E801F",
INIT_25 => X"A38BF8FC000000000000000000000000000000000000000000002ABEFAA80001",
INIT_26 => X"7155BC2A87092AAFA9257F1C5BC00AA5D7FF8EAA57803AEBAF7F5D74AAA2A03A",
INIT_27 => X"BFBC7EB8005B55A85B555EF095F50578085BE8FC7A3F00516DA2D5451D7EBDB4",
INIT_28 => X"0975FFAAA1521FF492BF8F40B6AAB84AF555168A00EA8000150A801C01C7142E",
INIT_29 => X"2EBAE28168ABAA2D43D568BC5400168E90E2F412BEAE3D542A004380124921D2",
INIT_2A => X"2FA3AA28EA8168A954100071D2E90A855C7A00A38F6DE05B40480557A95A3A1C",
INIT_2B => X"16D1EAE925EA0BFEBF4AA09217F490568417085147B50A80095178157FEFA074",
INIT_2C => X"000002D57AAA8402A8743DBD202DA95568A95E800A8F57F6DA971F8F7FFFA42D",
INIT_2D => X"AAFFD1564BA2282BFA02A2C28000000000000000000000000000000000000000",
INIT_2E => X"5EFA87F57555AAFBD7555FFAE95408A8FDC31AD017D34ABA5D7BEAAAAD786BCE",
INIT_2F => X"C2087383F79A5046A37B55F38415555797D63BFF007F8B2B2D97D483AFA7BD9F",
INIT_30 => X"42000D382964A92B401E71D7581C33172EC0A0300A6AEA8FAF0451CA001D4845",
INIT_31 => X"C8365A2FD5E04AA5780A8AAAD7AC3CA02003BEBBA7D7463CC508D07577BAFBD5",
INIT_32 => X"0621F562B1122DA70C3808458881056A5502AA150502828811FCD4EABDB1DFDF",
INIT_33 => X"96D55BBAAC55EAFAF86D35E4A92B4460D15060374FF72AAADF24559515705079",
INIT_34 => X"007FC0000007FC0000007FC07AAF12E00505D3FDF6A03D4BFB79AFA4C5CB5F58",
INIT_35 => X"0007FC0000007FC0000007FC0000007FC0000007FC0000007FC0000007FC0000",
INIT_36 => X"00000000000000000000000000000000000000007FC0000007FC0000007FC000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000040000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"CA1800080848B0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000010822C00803804000001999EF9C00040B0002000001000640200001018",
INIT_05 => X"0000400244000000014200004000000004000000001000032000200002100800",
INIT_06 => X"208500000080412804100CB08000302220080408010000202000000404100844",
INIT_07 => X"5AF6FEF002230018010860C1833C460044204C000008A0041000080008202800",
INIT_08 => X"8D22C0F55000010000524481890BC000263000188AAAA10F8C1830562B25FC4C",
INIT_09 => X"B102002E20013600022D8819000000A000110A4000002C204000240420001000",
INIT_0A => X"02605C1C1108481200C000002040040820000020104100028800002801041001",
INIT_0B => X"081001004010810510040802040102008100200800A1100707040101E20BE0B0",
INIT_0C => X"58000003C0F000A000C4000003C0F000A000C0000012187087010AE4B0000000",
INIT_0D => X"04000003C0F000A000C4000003C0F000A000CC4200002F08E03080000010F180",
INIT_0E => X"0000000AAC00680000001F10E038000000078808C00000023461C0E000000127",
INIT_0F => X"5200040A00D000000202090C281F201803000000240218C0044200001E187806",
INIT_10 => X"400012900001EC03F000000000392100B00048230C200009A000130320480002",
INIT_11 => X"308000000961002880204A901C0E00000002C9000260640900004D0000904618",
INIT_12 => X"5C0C0312A002000000083881002880025A0A3C020000002A8400B00007806070",
INIT_13 => X"04080830008010468220A00008D0000801046004308A18500002012800090428",
INIT_14 => X"0840280206089000004090110200000000001454000200828008081110084000",
INIT_15 => X"4191AC191AC191A4191A00C8560C8D2910000060901010401E13405111220000",
INIT_16 => X"0410028000100800140000002004103224002006406401918C191AC191A4191A",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200800041",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"0000000000000200802008020080200802008020080200802008020080200802",
INIT_1A => X"2431A589945201924924B060D757DF8A94102E038728287452B4008A04000000",
INIT_1B => X"75BADD6EAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8A28A28A28A28AB20",
INIT_1C => X"974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D6EB75BADD6EB",
INIT_1D => X"00000000000000000000000000000000000303FFFFFFFFFFFFFFC00000BA5D2E",
INIT_1E => X"FDFFFA2FFD74000855555FFFFFFC01FF087BE8BFF5D2AAAB5555554000000000",
INIT_1F => X"EBFF455D04175FF5D7FEAAAA002ABDEAA5D2EBFFEFA2D17DEBAF7D1574BAAAFB",
INIT_20 => X"8415400005540155F7D16AB45002EA8ABA005540145557BFDEAA5500154AAAAA",
INIT_21 => X"5003DE00A2FFFFFEFAAD57DE00082AAAA00082A820BAAAD540145F7D5574BAAA",
INIT_22 => X"F7D5554AA5D2ABDEBA082A821455D2EA8B455D2A975EFF7AEBFF550055555FF5",
INIT_23 => X"FFF84155FFFFFFFFF55AAAABFFFF5D556AB45A2D16AABAAAAEBFE10AAFBD7545",
INIT_24 => X"10FF84174BA552EBDEBA0004020AA5D04155FFAAFFEABEFA2FBEAB455D7BD55F",
INIT_25 => X"F47015A800000000000000000000000000000000000000000000175FFF7D1400",
INIT_26 => X"FEAAF7D5524AAA2F0BAF7FABDFC7E10005F525D74BFBC51FF1471E8BEF55242F",
INIT_27 => X"50492490E17EAAA2AAB8F4515043DFC75575C7000B6AEBAEAA5D2EBDFFFBED17",
INIT_28 => X"B6FB6DF7DFD5038ABA140A2D00554517DEBDB6FB55142A8708202FBD257F1C75",
INIT_29 => X"AABFF55BC5B555C74B8A38E38085BE8B47A3A00503D1420AD000B420820AAE2D",
INIT_2A => X"AABD21EF1C2FEA5FDEBDB505FA4920AFE10082E925555F8FFDE38087FC51C7F7",
INIT_2B => X"1EFBFDBFF5FF1C00BF5D25475C7B7FEAFF45BEAABA4AF555168B68FEDF6AB52A",
INIT_2C => X"00000151EAE3D542A004380124921D20BFFFA0AA17AEB8BFF155552B6F5E8BFF",
INIT_2D => X"FF55516ABEFDD003EFE5093DC000000000000000000000000000000000000000",
INIT_2E => X"2BA5D2ABDFFFF7D57DEAAFFD5420B2A2D37DB07A3D795000087BC01458AFBC11",
INIT_2F => X"D608897FD610D01151C610592A974BAFBAC28B55550434D555C53E0CE2AAA874",
INIT_30 => X"3FE102400144ABAAFFF7DE772FDD56588042F72EF0851575FFAAFBDD5542B2ED",
INIT_31 => X"F6A81A239501755F504BDF557D79431FD006EABA100F3D68FFFAABAC20EF0400",
INIT_32 => X"55EAF57FF957CAAA7FABF7DFD0C6A7DFFFA07FC04EA0006BFE007E2E8315DD02",
INIT_33 => X"FADF6900FFFF68BEFDFFB4B1FE5551141E78A02803158517BD745AEAEA8FAF0C",
INIT_34 => X"0000000000000000000000165BAFBD542000D382964A92B403EE18D5408A6F2A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000040000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0812",
INIT_01 => X"A145A00810790848048044A54E404340404000720885800802000906E4910200",
INIT_02 => X"5C010802020408040C455850AA055254090541A111200A104A0000000908B510",
INIT_03 => X"182002200C00004485264A001214912802150020218808002440854288890550",
INIT_04 => X"210302008014100120806B08702010102722C9E0412200651102418214049492",
INIT_05 => X"48416A98042912208552102442884882A58A08011290A1120A81230240018DCA",
INIT_06 => X"12800554528021C8023A28000031240048000100001170000155414109102066",
INIT_07 => X"000022104040810089080810211A04480420420154800088096A0EA8C0222080",
INIT_08 => X"080198C105424705510A08828A0B19080428040080A0A10F8102049300000804",
INIT_09 => X"3165541CD54822160A89E89020AA8AC4CA1D39CE215264B04040002400B80688",
INIT_0A => X"280201840548C80001C568146000001012D40D7182411080153801004800B057",
INIT_0B => X"4812050000080114100206000100818100900640C04C20104101021C00000310",
INIT_0C => X"00A00000010000A01001400000010000A0100801407234E34C1A980001552055",
INIT_0D => X"01400000010000A01000A00000010000A0100038000000000800000000405000",
INIT_0E => X"00000040A00002600000000010000000004608000850000000080000000001A0",
INIT_0F => X"400020C4000200420040000000001000000000002408000000A1000000020000",
INIT_10 => X"00001A04940000000000000020012800018000000000000D0288000000000003",
INIT_11 => X"0000000021480000508000000000000000400951000000000000681300000000",
INIT_12 => X"00000000000000000008600800004C000000000000000082A000015000000000",
INIT_13 => X"80004012C06000018004342AA000700000000000044000500000000022101800",
INIT_14 => X"958100134200904487400010022005E0110D524029263100009200151409130A",
INIT_15 => X"C9013C9011C90134901144801A4808AD4451394CD0391A541593C04B59084008",
INIT_16 => X"010400A0A890684444240120C0071420344423040240450114901149013C9011",
INIT_17 => X"080601806018060180200802008020080601806018060180200802048026C000",
INIT_18 => X"8000080001804018040180400800008000080601806018060180200802008020",
INIT_19 => X"1F83F03F03F00180401804018040080000800008000180401804018040080000",
INIT_1A => X"E90C042CB002102CB2CB2EE00271AE180616A85246C77250C7D00022012F81F8",
INIT_1B => X"28944A2504104104104104104104104104104104104104104104104104104608",
INIT_1C => X"128944A25128944A25128944A25128944A25128944A25128944A25128944A251",
INIT_1D => X"000000000000000000000000000000000003C3007FFFFFFFFFFFCE3F00944A25",
INIT_1E => X"EAA1055042AA105555421EFFFD568AAA002EBFEBA550002000AA800000000000",
INIT_1F => X"AA8BEFAAAE975FFA2D5555450851574000851554BAFFAE801FF087BE8BFF5D7B",
INIT_20 => X"2EA8AAA5D2EBFFFFA2D1554BAF7D17FEBAAAFFFDFFFA2D57DE10557BE8ABAF7A",
INIT_21 => X"D04175FFFFD5574AAAAAA974BA082EA8BEFAAD555555F7D568ABAF7D5574BA55",
INIT_22 => X"085557410F7AA97410087BD55FF087FEAA10A2FFEAAAA552AAAAAAAAAABFF455",
INIT_23 => X"05D7FE8B45F7FBFDE00085540155F7D56AA00007FEAA000055401555D7BFFE10",
INIT_24 => X"00082A820BAAAD540145F7D557410AA8428A10550017400550402155A2803FE0",
INIT_25 => X"000E28A80000000000000000000000000000000000000000000017400082AAAA",
INIT_26 => X"01FF1471E8BEF5574AFA00010ABFA38555F401D74BD16FAAA002ABFEAA550E82",
INIT_27 => X"FF400417FEF082F7AAA8BEFE2AA955EFA2DB5757FEAFBD2410005F57482E3AA8",
INIT_28 => X"F6DA82F7DF520385D2FE80AA5D2EBDFD7BED1574AAF7D5524AAA2F1FAF7FABFB",
INIT_29 => X"24ADAAAB6AAB8F455784155C75575C7000B6AE95492082EADBFFBEDB55555E3D",
INIT_2A => X"051C05571474024A81C5557578EBA087400007FC21C7005B6FB47F7A438E925D",
INIT_2B => X"E10A001FFB40038F68F7F578F7FFEF568E2808554717DEBDB6FA3D0075EDA800",
INIT_2C => X"000001043D1420AD000B420820AAE2DB4716DF7DFFDE381D716FA15550015428",
INIT_2D => X"AA002ABDEAA552A80010AAA88000000000000000000000000000000000000000",
INIT_2E => X"800087BD5410AAAA801FF55556ABEF5D517EEE00828FDEBA5D7BC015582D57DE",
INIT_2F => X"A2B2A3D169B07A3D7BFE10597BFDE00AEAC28BFFAAAE955EFAAFBC15F5A3D7D6",
INIT_30 => X"BDFEFFFFBC1154AAFFFFE107FF9D72A20842080BA5D2ABDF55F7D575EAAFFD50",
INIT_31 => X"97CF4780286A2105D2A3FEBAFFAC28B555504145555A53C00B2A2AA02000082A",
INIT_32 => X"FFFDA02003FFDEAA8557D65550915544AA5D51574EAA28015400547FC315D007",
INIT_33 => X"16F9E2555500174AA282E20BFFFF842AAAAADD5699ADABD5A8AAA0051575FFA2",
INIT_34 => X"0000000000000000000000030EF04003FE102400144ABAAFFD75E7F2BDDD2B80",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000080000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380202",
INIT_01 => X"200C9A424080216D3C2462C99E104B49404040028804A0080A000416A8D90A0C",
INIT_02 => X"4809A902031800444461089C66E331352180D468B8240E600C0081110B80ACD0",
INIT_03 => X"DA16C2210C0001D231A30A0648C68428320066010A80881068A80C401CC46330",
INIT_04 => X"2088601DA82700EC92307064A3756910088469A01C250210990240420E005A48",
INIT_05 => X"2D2060182414411A314A0A02C18C01B9854368080A506912018C2502484038D1",
INIT_06 => X"16801CCCAA8061E8061C0D008020140520080769000420202133CCC50C110804",
INIT_07 => X"5800B65040630008810C20508138071604A461833280038C89904E6400232008",
INIT_08 => X"0800906010521D1CC80204918949540C061000088000A90F840A50963A017845",
INIT_09 => X"A037A02C68552A35620C88900A69876100810A6A84C82C400040300D40D20A48",
INIT_0A => X"062A10B40042C80000CCE4CC2045051913208CE80243048008204100402079CC",
INIT_0B => X"C81301004C18912102060C0207010201C190200400A401042D00F15884030170",
INIT_0C => X"0190148000000800100450148000000800100401CB33494594532980733322CC",
INIT_0D => X"05101480000008001004F014800000080010051C000040000000000000480000",
INIT_0E => X"00000044000001680180400000000000014000000B1004090000000000040080",
INIT_0F => X"00812E44000024400140800280000000000002000008000001B0000040000000",
INIT_10 => X"0002080CCC0002000000000020401000034010480000010402D8040440000041",
INIT_11 => X"00000000601000064180104400000000004100570080880000082015C0209000",
INIT_12 => X"00820080000000000100401000061C0001000000000000904000094C00201800",
INIT_13 => X"4408400000A26285A03224E670094008010000004444010E2050000420801880",
INIT_14 => X"4DC10283429294408740C0B48202854C011CD75C0102A30400A8891451284B26",
INIT_15 => X"4901A4901849018C901A648056480C2D4449116DC0115C41159B655F112AC008",
INIT_16 => X"0510000000DA690C1D20030BA0011421B404220402404501A49018490184901A",
INIT_17 => X"280803808038080380803808038080380C0280C0280C0280C0280C0680C28051",
INIT_18 => X"00C0280E030080380A030080380A030080380C0280C0280C0280C0280C0280C0",
INIT_19 => X"B556AA9556AA830080380A030080380A030080380A0200C0280E0200C0280E02",
INIT_1A => X"742C000A981E80249249206018F18E0C85142822266800586291000A844D54AA",
INIT_1B => X"A9D4EA7524924924924924924924924924924924924924904104104104104A20",
INIT_1C => X"1A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A753A9D4EA753",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF849010D46A35",
INIT_1E => X"42000AA802AA10F7D57FEAA557BE8B45A2D5555EFAA800015508000000000000",
INIT_1F => X"BC0155A280021EFA2FFE8B4555042AA105555421EFFFD568AAA002EBFEBA5551",
INIT_20 => X"D5574000851554AAFFAE801FF087BC01FF5D7FEAA10550402000AAD56AAAA557",
INIT_21 => X"AAE975FF005540145A2D157410AAD17DFFF5D0400010AA842AAAAFFD542000FF",
INIT_22 => X"F7AE975FF080428B455D7FFDEAA5D55574BA00517DE105551420BAF7AAA8BEFA",
INIT_23 => X"F007FFFEAAAAD5554AA552EBFFFFA2D5554BAF7803DEBAAAFFFDFEFAAD57DEAA",
INIT_24 => X"EFAAD555555F7D568ABAF7D5574BA552E800BAAAAE800AA087BD5555552A821E",
INIT_25 => X"155080E800000000000000000000000000000000000000000000020BA082EA8B",
INIT_26 => X"FAAA002ABFEAA555E02000E28AA8A38EBD578E82E975EAB6DBEDF575FFAA8E02",
INIT_27 => X"87A38AAD56DA824975C217DAA84021FFAAF5EAB55EBAEADA38555F451D7EBD16",
INIT_28 => X"E2DABAFFDB47412ABFE90410005F57482E3AA801FF1471E8BEF5575EFA00012A",
INIT_29 => X"5F47082E3AAA8BEFA02A955EFA2DB5757FEAFBD2400BED57FFD7410E05038BE8",
INIT_2A => X"2F1FAF7FABFBEAE2AEBA4974871C043AB6D4975FFEBA5D71D742A407FFFE0055",
INIT_2B => X"1C75D25C74920821D708757AE2AA3FFC04AA552EBFFD7BED157482F7803AEAAA",
INIT_2C => X"0000007092082EADBFFBEDB55555E3DF6DA82F7DF7AE38497FC00BAB6A485082",
INIT_2D => X"FFFFFFD75FFAAAE8014500288000000000000000000000000000000000000000",
INIT_2E => X"EBA5D7BD5545A2D57DEAA002EBDEAA557BC0010AAA8A8ABAAAD568A1020516AB",
INIT_2F => X"29EF5C517EEE00828D74AAFBD57DE000057C21FFAA80001FFAAD57EB55A2A8AB",
INIT_30 => X"7DF55082E974AAFFAABDEBA77FDD66A0ABBDC2000087BD5410AAAA801FF55556",
INIT_31 => X"7C14100957FF6105D7BD5400AAAC28BFFAAAE955EFA8FBC15E5A3D5D7400FFD5",
INIT_32 => X"D1554A8FFC42AA10A7D169F57ABD7FEEBAAA841550555002ABFF54517EEB25D5",
INIT_33 => X"96F014AAFF84154105555C215500000014558557FA42A3D7020BA5D2ABDF55F7",
INIT_34 => X"000000000000000000000015400082ABDFEFFFFBC1154AAFFFFE10FFF9DF2020",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000040000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204002",
INIT_01 => X"010398000008004C1C20650E1E104348403008418984014902030006A0910200",
INIT_02 => X"480108A200000000444048E41E80F00A4104311868200200080000000988A390",
INIT_03 => X"0CA08220080000D004060A0240101028270012603000000030808C0208C000F0",
INIT_04 => X"4403A609A055306BC2C0735810CEE5100A0A40E06B8360E3808241D03845D002",
INIT_05 => X"ECE0498800791403AD3038AE079059A790E245819A41E4120BAB87800001D312",
INIT_06 => X"06000C3D220003E0001A210088B1008C4004034912120000010FC3C00000A064",
INIT_07 => X"5000220440000000090800002118400204206100F040018019004B8001232088",
INIT_08 => X"0810884441123323C0424180880B0108002000000880890F9000041200000845",
INIT_09 => X"230B6715A4786E0F5A8C889031EF9F45D884794FA03A24781840100D000E1140",
INIT_0A => X"0C4202200142400004DC3C82600401003200872003FB1400082840001022003C",
INIT_0B => X"C800940008088034040000010000808140901000C00001008800A01814000840",
INIT_0C => X"02E0100000000800000620100000000800000001C07261841840310240F070C3",
INIT_0D => X"0680100000000800000760100000000800000435100040000000000000080000",
INIT_0E => X"00000004000000D8008000000000000001000000155000080000000000040000",
INIT_0F => X"000100EC00004002214000008000000000000200000000000094100040000000",
INIT_10 => X"000200010C000200000000000040080005800008000001000368000040000040",
INIT_11 => X"000000004008000448000040000000000001007C000008000008001D00001000",
INIT_12 => X"000000800000000001000008000017000100000000000010200002C800000800",
INIT_13 => X"0000549000027200800E271E00288400800208004804C0080000000052800800",
INIT_14 => X"454000924280D144B14041340A880EC51160525C0022510006BE1002C6150F5E",
INIT_15 => X"010C1010C1010C3010C14086980861AD447F2201D899BA403593514B59A30088",
INIT_16 => X"010448002098694C15204369E00116203445E3443043410C5010C3010C1010C3",
INIT_17 => X"180000006018000000200804010020080400002018040000600800010064E000",
INIT_18 => X"8060000001000008060180201000000040180001006008000100201804000020",
INIT_19 => X"934D964C32698000401802008060000401000008060080201004000000080201",
INIT_1A => X"0991A185145019A28A289830C700FC0A0002870BB5ED0B34504048828464B261",
INIT_1B => X"351A8D46AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8A28A28A28A28AF4C",
INIT_1C => X"8341A0D068341A0D068341A0D068341A0D068341A0D068341A0D46A351A8D46A",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8EE3EC1A0D06",
INIT_1E => X"40155080000155FF843FFEFAA84001FF5D043FEAA5D55420AA002A8000000000",
INIT_1F => X"A80010FFAE975FFAA80001EFA2AAAAA10F7D57FEAA557BE8B45A2D5555EFAAD1",
INIT_20 => X"AAAAA105555421EFFFD568AAA002EBFEBA555542000AA80001555D04174AA002",
INIT_21 => X"280021EFA2FFE8B45F78400145FF842AAAAA2AA800BA5D51555EF002AA8BFFAA",
INIT_22 => X"00003DFEF080428B455D002AABA5D2AAAAAA5D2E82000AAD568AAA557BC0155A",
INIT_23 => X"FAAAAA8BEF552E820000851554AAFFAA801FF087BC01FF5D7FEAA105D0428B45",
INIT_24 => X"FF5D0400010AA842AAAAFFD542000FFD57DF55A280154BAA2FBE8AAAF7AA821E",
INIT_25 => X"092142E00000000000000000000000000000000000000000000015410AAD17DF",
INIT_26 => X"AB6DBEDF575FFAADE02155080E85145E3803FFEFA284051D755003DE92415F42",
INIT_27 => X"851455D0A124BA002080010FFA4955C7BE8E021C71C0A28A38EBD57DE824975E",
INIT_28 => X"B505D71424AABD7F68E2FA38555F451D7EBD16FAAA002ABFEAA555F42000E2AA",
INIT_29 => X"D56DA824975C217DAA84021FFAAF5EAB55EBAE82145F7802AABAA2A480092415",
INIT_2A => X"575EFA00012ABFB6D080A3AFEF080A2FB45490E2AA824924AAA92550A07038BE",
INIT_2B => X"AAFFEAA00F7AE821D7B6A02FBC71D0E10010005F55482E3AA801FF1471C01EF5",
INIT_2C => X"0000010400BED57FFD7410E05038BE8E2DABAFFDB6FA12ABAEBDF7DAA80104BA",
INIT_2D => X"4555043FE10087BC2000552C8000000000000000000000000000000000000000",
INIT_2E => X"ABAAAD57DE1000516ABFFFFFBD75FFAAFFC0145002897555A2803FFFFAA84175",
INIT_2F => X"DEAA557BC0010AAA895555042E820BA080400010FF8017545F7AE821455D2CAA",
INIT_30 => X"2AAAAAA8002010007FC0155D5022A955FFACBFEBA5D7BD5545A2D57DEAA002EB",
INIT_31 => X"43CAB0552C97CAAFFD57DE000057C21FFAA80001FFAAD57EB55A2A880155F780",
INIT_32 => X"AA801FF5555421EF58517EAB00028A9BEF002EAABEF002EBDF45542AAAA00080",
INIT_33 => X"A90FDFEFA280020BAA2FFEAA10FFAE82145F7803CFE55D2CC2000087BD5410AA",
INIT_34 => X"000000000000000000000002000FFD57DF55082E974AAFFAABDEBAF7FDDE6A0A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000080000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A337A20E07C0C1E006",
INIT_01 => X"295FBC448000804C5C6A60000C34C26841280A00084000C8C212802EE2953235",
INIT_02 => X"C809AD5EB118E640A4D158FC011FF0002080000082E8C66609DB7DDDCB1FA036",
INIT_03 => X"4A120E4C3A4C90D214A35E824852857A0A20640A88800000B8E0FC52A884500E",
INIT_04 => X"001440809A2604005934800041110A71E290E8B010DB221C662AE22DC0AA3448",
INIT_05 => X"12026A2A1B88C31841CDC451B860A6507BEBD18A65AE10571450DE8112522449",
INIT_06 => X"80752C03736281D628398CD0A4C894EA2054237F271331095100D82D0C2C82A2",
INIT_07 => X"5E64B66BD6231CC81529A356AD3AC601C57FF54FF149A46490261C4B39203F70",
INIT_08 => X"AD0099410015814FC602C4B1B93947F8621030C800001D7FA46A95172E937835",
INIT_09 => X"2C836D35B68D26C082DE9AB88C104020000208401807B78739010C04E17F5014",
INIT_0A => X"082099129008F25615C3FC01A2102109204C28B6706168128920C469E7C00A00",
INIT_0B => X"E92C23E210A0B246C2234010A108D0042811461C0401502644A40106C14FD22A",
INIT_0C => X"E00BF1BFE1F000BE1FC40BF1BFE1F000BE1FC80028120800800100653FF0313F",
INIT_0D => X"040BF53FE1F000BE1FC40BF53FE1F000BE1FCC806FFFEF0AE83080E2AEF2F1F1",
INIT_0E => X"013879FAAF8FC003FEDF5F12F0380231F0FF963F00A7FBDF3669C0E008C3CBFF",
INIT_0F => X"F2008022CBAC8B9DDEB779BEA91F30180309A0F83FEAB8FC7C006FFFDF1A7806",
INIT_10 => X"4131BF940DFFFE03F00003F03FB929E9C19BE8EB0C2098DFE2EF7B2760483137",
INIT_11 => X"3080E29F3B69E9F4427EEED41C0E004C72FEC95DEFE46C090626FF1537F15618",
INIT_12 => X"FC0E0392A0024B83F07F7989E9F01DFFFB0A3C0202B877EAA7A7C1CBFFD07870",
INIT_13 => X"C0404020040001C4E7F1787E0C8028514885C566241902508C83A7D1B7EFAC6D",
INIT_14 => X"4DF46A170F92C7E20F0430938008AC38C4184B100136858C9298A8560688F4C1",
INIT_15 => X"6B8C86B8CE6B8CA6B8CC15C6435C670C10EB4124D2B3903BF5C9710C1191DCA0",
INIT_16 => X"2030461200984D041C40208400230E71B3104E5636E3178C86B8CC6B8CA6B8CE",
INIT_17 => X"0040118401184610042110401184410846110421104010844118421504238200",
INIT_18 => X"8441184011844100461004211046100461084211042100441084011842100461",
INIT_19 => X"DA6924965B4D1004610840118401084410840110421004610046110421084410",
INIT_1A => X"FF9FBFAF2DDA3B9E79E7BED9CFEF73B6FFE74FC3F78FFF6DB7ED438A183124B2",
INIT_1B => X"DDEEF77BBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEDFD",
INIT_1C => X"BDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BB",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF853FB5EEF77B",
INIT_1E => X"020AA002AAAABA555140155087FFFFEF00042AB555D2E955FFF7FFC000000000",
INIT_1F => X"E975FF5D5568B555D7BD5545FFD540155FF843FFEFAA84001FF5D043FEAA5D04",
INIT_20 => X"FFEAA10F7D57FEAA557BE8B45A2D5555EFAAD5401550800001FF5D00001555D2",
INIT_21 => X"FAE975FFAA80001EF002AAAABAF7D168A10A2D17FF45A2FFC0000AAAE974AAFF",
INIT_22 => X"F7803DF55FFAEBFE005D2EAAB45557BD55555555401555D04174AA002A80010F",
INIT_23 => X"5552E955EF5D7FEAA105555421EFFFD568AAA002EBFEBA555542000A28028BFF",
INIT_24 => X"AAA2AA800BA5D51555EF002AA8BFFAAAA820AA5D517DF55082E974BA087FE8B5",
INIT_25 => X"5C7F7FBC0000000000000000000000000000000000000000000000145FF842AA",
INIT_26 => X"51D755003DE92410F42092142E28ABA5D5B4516D007FFFFFF1C042FB7D492A95",
INIT_27 => X"851C75D0E02145492E955C75D5F6DB55497BD5545E3DB45145E3803AFEFA2840",
INIT_28 => X"BC7028A2AA95492FFFFE8A38EBD57DE824975EAB6DBEDF575FFAADF42155082E",
INIT_29 => X"0A124BA002080010FFA4955C7BE8E021C71C0A2DABAF7D16DA28A2DB7AF7DB6F",
INIT_2A => X"55F42000E2AAA8BEFE3843AF55E3AABFE105520AFB45557BD5555415F4514549",
INIT_2B => X"082E954AA087FEDB7D5D2A155D7157BEFA38555F451D7EBD16FAAA002ABFEAA5",
INIT_2C => X"0000002145F7802AABAA2A480092415B505D71424821D7F68E07082495B7FF7D",
INIT_2D => X"EF5D003DFEF002E95555F7FDC000000000000000000000000000000000000000",
INIT_2E => X"555A2802ABFFAA841754555043FE10082A82000552CAAAAA5D7FD75EF087BFDF",
INIT_2F => X"75FFAAFFC0145002895545552E80145002E955455D7BFDF45007FD7555A2F9D5",
INIT_30 => X"7FEAAAAFFEABFFF7FFD54BAA2AA95410F7FDEAABAAAD57DE1000516ABFFFFFBD",
INIT_31 => X"BD55550879D5555002E820BA080400010FF8017545F7AE821455D2CBFEAAFFD1",
INIT_32 => X"D57DEAA002EBDEAA557BC0000AAA8A8BEFA28028B45AAAABFE0009043FF555D7",
INIT_33 => X"FAC97400087FFFFFF002E954AA087BFFFFF5D2E975455D7DFFEBA5D7BD5545A2",
INIT_34 => X"000000000000000000000000155F7802AAAAAA8002010007FC0155550222955F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000300000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B0061A258A2840112C03002C180004003220200403302301C0381A0082",
INIT_01 => X"860041C838394848008100000042026041000000090800090210010000510204",
INIT_02 => X"080108220C1000004464080000C008010000000001243240080080000988A050",
INIT_03 => X"080000010C23404080020A600200002983800504488000103080050C08C10000",
INIT_04 => X"0040504280A682104011230010000010002040E9102050101000400A00003000",
INIT_05 => X"0409400984008000414A00014000002004100020005004020010204044802800",
INIT_06 => X"301223FC028911E8911900000224200248A653E908C0248489FF000809108000",
INIT_07 => X"0000220441820000090C080001184400142040200E824008900008000220600A",
INIT_08 => X"1A18946451007FA0380200808809010C182000000000090F8100001220000804",
INIT_09 => X"300240B4A409223F020988100808200490142B441BF82C20401481540A000008",
INIT_0A => X"264285180542408000D001BE090693912000002004410489080001100017E2FD",
INIT_0B => X"091081090A4491A40052A129519428CA142288010A5A21214601F01A220602A0",
INIT_0C => X"18100400000000A00034100400000000A00033A00813004104020818800F2400",
INIT_0D => X"F4100080000000A00034100080000000A0003142000000000000000000055D00",
INIT_0E => X"00000001E8002900010000000000000000066000C20004000000000000000120",
INIT_0F => X"4D240C2000502000000080000000000000000000240146800142000000000000",
INIT_10 => X"00001260F0000000000000000007F00032201000000000091A00040000000002",
INIT_11 => X"0000000005D00008958010000000000000003F4000008000000048D240008000",
INIT_12 => X"008000000000000000082670000CC0000000000000000007C000301400200000",
INIT_13 => X"0120849A5250101482202301F05101202420000810C219500150002800101280",
INIT_14 => X"454110030212C140011204D020880C000018431DE802015022A62A1596C8B580",
INIT_15 => X"016C2016C2016C6016C440B6000B600C446B0104D09192013589701C59800002",
INIT_16 => X"51804A0028904C425016040820978221B0000005B05B416C0016C0016C4016C4",
INIT_17 => X"8CA3294A528CA328CA1294A528CA3284A5294A728CA3284A529CA728CA100508",
INIT_18 => X"CA3284A129CA7294A328CA1294A729CA128CA329CA5294A128CA3294A5294A32",
INIT_19 => X"1C71C718638E28CA529CA7284A128CA7294A528CA1284A729CA1284A3284A529",
INIT_1A => X"ED9DBDAFBC5E9BBEFBEFBEF9CFF1FE1E9F52AFF9F3E77B7CF7F40A00107638C3",
INIT_1B => X"FCFE7F3F8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E76C",
INIT_1C => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9",
INIT_1D => X"00000000000000000000000000000000000303007FFFFFFFFFFFC61AC8FE7F3F",
INIT_1E => X"955FFF7FFC21EFF7D17DEAA5D2AAAAAA5D557DE105D2EBDF55557FC000000000",
INIT_1F => X"03DEAA5D5568BEF5D042AA10A2AAAAABA555140155087FFFFEF00042AB555D2E",
INIT_20 => X"5540155FF843FFEFAA84001FF5D043FEAA5D00020AA002A82145555542010FF8",
INIT_21 => X"D5568B555D7BD5545FFD568AAA5D00154AAAAD1420BA00557DF455D7BFFEAA55",
INIT_22 => X"F7843FF55007FFDEAAA284020BAAAD168BFF0800001FF5D00001555D2E975FF5",
INIT_23 => X"5AAAEBFE10FFFFEAA10F7D57FEAA557BE8B45A2D5555EFAAD540155080000000",
INIT_24 => X"10A2D17FF45A2FFC0000AAAE974AAFFFFC21EF5551401EFF7842AA00FF841754",
INIT_25 => X"F45497FC000000000000000000000000000000000000000000002AABAF7D168A",
INIT_26 => X"FFFF1C042FB7D492A955C7F7FBC71EFFFD57FE825520ADA92495B7AE10412EBF",
INIT_27 => X"0716D415F47000F78A3DE92415F6ABD7490A28A10AAAAA8ABA5D5B4516D007FF",
INIT_28 => X"F78F7D497FFFE925D5B45145E3803AFEFA284051D755003DE92410E02092140E",
INIT_29 => X"0E02145492E955C75D5F6DB55497BD5545E3DB6AA92550A104AABED1470AA005",
INIT_2A => X"ADF42155082E87038FF8038F6D1C7BF8EAAAA80020BAA2DB68BC7140E051C75D",
INIT_2B => X"FF8428A00E38412545AAAE3FE10A3FBE8A38EBD57DE824975EAB6DBEDF575FFA",
INIT_2C => X"000002DABAF7D16DA28A2DB7AF7DB6FBC7028A2AA95492FFFFC71EF415F471C7",
INIT_2D => X"00007FEAA10002ABFF450079C000000000000000000000000000000000000000",
INIT_2E => X"AAA5D7FD75EF087BFDFEF5D003DFEF002E95555F7FDD55EFF7D57DE005D003DE",
INIT_2F => X"FE10082A82000552C955FF007BD5410FFAABFE00087BE8B45082EAAA10A2A8AA",
INIT_30 => X"820AAF7D5574AA087BEABEF007FFDE00557DD5555A2802ABFFAA841754555043",
INIT_31 => X"BEAB55552C95545552E80145002E955455D7BFDF45007FD7555A2F9EAA005D2A",
INIT_32 => X"516ABFFFFFBD75FFAAFFC01450028974BAFF842ABFF557BE8ABAA284020BAA2F",
INIT_33 => X"7FDD55EF007BD5555F7802AA10AA8000145AAAEBFE10A2F9EAABAAAD57DE1000",
INIT_34 => X"00000000000000000000003FEAAFFD17FEAAAAFFEABFFF7FFD54BAA2AA95410F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000240000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C024504188000003000000003302300C018180006",
INIT_01 => X"020008422008604D042080000211024840000000080000080200080000110204",
INIT_02 => X"4801082048100000444008040080000041000000000222400800000009000010",
INIT_03 => X"0802030288A148D0000208424000002103006400088000003080000408C10000",
INIT_04 => X"00004000890600004032030010000010008060E4100000140006500800403040",
INIT_05 => X"0400400080000018414800810000002000000000004000328010000080882000",
INIT_06 => X"281A8001220021E0021803000224200200000360888420000000100808000000",
INIT_07 => X"5000220409020000090800000118040014A061200052500810000C490323208E",
INIT_08 => X"1A9098411110014000424090980B0002102000000000010F8000001220000805",
INIT_09 => X"31024034A4092200820D899408000004D0143B4410002C800080020450800001",
INIT_0A => X"24028011444240A88CC00100200D0010200008B2066397014800221400140C01",
INIT_0B => X"080001000C008124000000000100008000100404204C25200451A01A00A620A5",
INIT_0C => X"1C0014800000F001E02C0014800000F001E021141213000000000010B0001000",
INIT_0D => X"CC0014800000F001E02C0014800000F001E022420000400004C3201C51040908",
INIT_0E => X"60078601084038000180400002C0E00E0E004100E000040900000B0380383400",
INIT_0F => X"08146800105100000000800284004160C0301D07001504820242000040000198",
INIT_10 => X"908C404AFC000200030F000FC00610103BE0104810C8462014F8040446120C88",
INIT_11 => X"C3201C608410100FD5801044013098038D00309F008088C2419100A7C0209021",
INIT_12 => X"00B2048902C0807C0E008450100FDD000100411C8107880440403DDC00201804",
INIT_13 => X"00100496406010A0A2002200125140000000221110C018066250402E32901A80",
INIT_14 => X"454214028220141530400910CA800900326790500002001444001C0050140A00",
INIT_15 => X"5120551205512055120708901A8901A104804000801212541403C15178008010",
INIT_16 => X"01004200A09A49445420000DC000152804C9A384814809201512015120151201",
INIT_17 => X"0004000000080200806008020000000000000020080200802000000000008000",
INIT_18 => X"0000000000802008000000000002008020000400000000000080600802008000",
INIT_19 => X"0002082080000100000802008020100000000008020180000000000020180200",
INIT_1A => X"0000000000000000000000000000000000000000000000000005428A14584104",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8DD9EC000000",
INIT_1E => X"BDF55557FFDE00557BEAABAA2AEAABEFF78015555AA801741055554000000000",
INIT_1F => X"BEAAAAAAD157555AA803FEBA5555421EFF7D17DEAA5D2AAAAAA5D557DE105D2E",
INIT_20 => X"802AABA555140155087FFFFEF00042AB555D2E955FFF7FFD5555557BEABFFF7F",
INIT_21 => X"D5568BEF5D042AA10A2AA955EFF7FFD5400F7FFFDFEFAA80000BAAAAA820BAA2",
INIT_22 => X"5D7FE8A000004154BAF780001EFAAAAA8B45000002145555542010FF803DEAA5",
INIT_23 => X"5AAD5555EF557FC0155FF843FFEFAA84001FF5D043FEAA5D00020AA002ABDEBA",
INIT_24 => X"AAAAD1420BA00557DF455D7BFFEAA5555575455D2AAABFF5551421FFAAD15754",
INIT_25 => X"4385D5540000000000000000000000000000000000000000000028AAA5D00154",
INIT_26 => X"DA92495B7AE10412EBFF45497FFFE385D71E8AAAAAA0A8BC7EB8417555AA8410",
INIT_27 => X"D056D5D75EABC7FFF5EAAAABEDF5257DAA8438EBA4155471EFFFD57FE825520A",
INIT_28 => X"0070BAA2A0870BAAA8028ABA5D5B4516D007FFFFFF1C042FB7D492A955C7F7FB",
INIT_29 => X"5F47000F78A3DE92415F6ABD7490A28A10AAAA925EFEBFFD2400EBFBFAFEFAA8",
INIT_2A => X"10E02092140E3DE924171E8A281C0E10482F784001D7AAA0AFB6D1C040716D41",
INIT_2B => X"4955421EFA2DF5557DAAD5D05EF0175C5145E3803AFEFA284051D755003DE924",
INIT_2C => X"000002AA92550A104AABED1470AA005F78F7D497FFFE925D5B525454124AFBC7",
INIT_2D => X"55A28015545A284000BA5D534000000000000000000000000000000000000000",
INIT_2E => X"5EFF7D57DE005D003DE00007FEAA10002ABFF450079FFEAA5D5568ABAA2842AB",
INIT_2F => X"DFEF002E95555F7FDC01EF55556AB55F7D56AABAF7FBC01EFA2842AABA085755",
INIT_30 => X"C2000A2FFEABFFAA84174BAAA80174AAAA862AAAA5D7FD75EF087BFDFEF5D003",
INIT_31 => X"43DFEF5D02155FF007BD5410FFAABFE00087BE8B45082EAAA10A2A8801FFA2FF",
INIT_32 => X"841754555043FE10082A82000552CBFE10085168AAA552A80010F78000145AA8",
INIT_33 => X"57DC014500003FF450051401FFA2FBD55EFAAD5421FF085755555A2802ABFFAA",
INIT_34 => X"00000000000000000000002AA005D2A820AAF7D5574AA087BEABEF007FFDE005",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0000040042840002C00000018000002700500030B3132000400812082",
INIT_01 => X"A14008420008204D042100000212026840000000180800080200090048510200",
INIT_02 => X"080108020090000004655C000080000051000000002402400800000009008010",
INIT_03 => X"0002000100300C408422420002108108028065044880001030808D4288C10000",
INIT_04 => X"0002504688A28210003100000000001002A0E88910A032541000090A00643040",
INIT_05 => X"04092A081400D118410A002140004020140001A9005000004810A1C0044D2800",
INIT_06 => X"0010EFFD228931C8931820002080258A48A653E00213248C98FFC0094910A222",
INIT_07 => X"4000220440120000090C0810210A040034A040000046180810000C4907036008",
INIT_08 => X"50D88C2450000140004200808809000C012000000000010F8102041320000000",
INIT_09 => X"2002002020010200828C88020800200040801A40100228A1585481544A804040",
INIT_0A => X"A20804802400C80080D0010029069290200008B20E2304086800400640200801",
INIT_0B => X"091084090A4C81240251A328D094684B34A288050A5828012009504420102180",
INIT_0C => X"080004801E0FF00010000004801E0FF000100220021200000000000080001000",
INIT_0D => X"000004801E0FF00010000004801E0FF000100440000000F517CF600000400104",
INIT_0E => X"E000004008100800010040ED0FC7E000004008804000040109963F1F80000080",
INIT_0F => X"0020040020100000000882431660CFE7C0F00000000800810040000000E587F9",
INIT_10 => X"B0000808000001F80FFF0000200008021040134473D800040010045C1F360001",
INIT_11 => X"CF600000200802028001102EA3F1F80000400002008B83D6C0002000802688E7",
INIT_12 => X"03F2DC2D1FC18000000040080202800004D5C3FD80000080200818000027928F",
INIT_13 => X"0122C01A52501094222002000110012064200008848218002100100C00004112",
INIT_14 => X"4500048240C08400841204D0A00089000100001DE9248104300294428148A480",
INIT_15 => X"4800048000480004800004002240020850884000901210140011C010312B888A",
INIT_16 => X"51A4C000889A4D0E1D7624086491800420044240020004004480004800048000",
INIT_17 => X"84A1284A128CA328CA328CA328CA328CA328CA1284A1284A1284A12C4A14E508",
INIT_18 => X"CA328CA3284A1284A1284A1284A328CA328CA328CA328CA3284A1284A1284A12",
INIT_19 => X"000000000000284A128CA328CA328CA328CA3284A1284A1284A1284A328CA328",
INIT_1A => X"4799B1A014503EB65B6594F14A87D78AF421448BB528AF75D640088884400000",
INIT_1B => X"7C3E1F0F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79EDFC",
INIT_1C => X"87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F0F87C3E1F0F8",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF834FA53E1F4F",
INIT_1E => X"174105555420000000021EFAA843DE00F7803FEBAFFFFC2000557FC000000000",
INIT_1F => X"43DE005504175FF08514014555557DE00557BEAABAA2AEAABEFF78015555AA80",
INIT_20 => X"7FC21EFF7D17DEAA5D2AAAAAA5D557DE105D2EBDF55557FD54AAA2AA955FF000",
INIT_21 => X"AD157555AA803FEBA55556ABFFA280154BAFF803DF45FFD17DFFFFFD56AA0055",
INIT_22 => X"002AAAAAAA2D57DF450004154BA087BEAAAAF7D555555557BEABFFF7FBEAAAAA",
INIT_23 => X"5FFD1555EFA2802AABA555140155087FFFFEF00042AB555D2E955FFF7FFD5410",
INIT_24 => X"00F7FFFDFEFAA80000BAAAAA820BAA280000AAA2843DE1008556AA00A28028B5",
INIT_25 => X"0285D75C00000000000000000000000000000000000000000000155EFF7FFD54",
INIT_26 => X"8BC7EB8417555AA84104385D5542038000A001C7A2803AE38FF843DEBAEBFFC2",
INIT_27 => X"D24BAA2AA955C708003FE285D00155FF0055451555D5F7FE385D71E8AAAAAA0A",
INIT_28 => X"B78FFFE3DF6DA284175C71EFFFD57FE825520ADA92495B7AE10412EBFF45497F",
INIT_29 => X"75EABC7FFF5EAAAABEDF5257DAA8438EBA415568BEFA28E124AAF7843AF7DEBD",
INIT_2A => X"92A955C7F7FBD54380020ADA82BED57DF450804104920875EAA82F7DB5056D5D",
INIT_2B => X"005F68A10BE802DB55E3DB555FFF68028ABA5D5B4516D007FFFFFF1C042FB7D4",
INIT_2C => X"00000125EFEBFFD2400EBFBFAFEFAA80070BAA2A0870BAAA80070BAA2803DE00",
INIT_2D => X"AAFF803DEBAAAFBC20BA55514000000000000000000000000000000000000000",
INIT_2E => X"EAA5D5568ABAA2842AB55A28015545A284000BA5D53420BA082E82155AA802AA",
INIT_2F => X"AA10002ABFF450079C20BAAAAE9754500043DEBA5D04175EF0855575455D7BFF",
INIT_30 => X"820AAFF802ABEFAAFFEABEFAAFFFDEAA0051555EFF7D57DE005D003DE00007FE",
INIT_31 => X"16AA10FFFFC01EF55556AB55F7D56AABAF7FBC01EFA2842AABA085768BFFA2AE",
INIT_32 => X"7BFDFEF5D003DFEF002E95555F7FDD74BA08043DE10F7D17FF55000000010085",
INIT_33 => X"A86174AAAA843DE00087FE8A00F7843FF45AAFFD75EFF7842AAAA5D7FD75EF08",
INIT_34 => X"0000000000000000000000001FFA2FFC2000A2FFEABFFAA84174BAAA80174AAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000100000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000006",
INIT_01 => X"000009801830084C182060000C104268413C0A61590001D90213C00000110200",
INIT_02 => X"680108200010000054400C000080000041000000010002400800800009082011",
INIT_03 => X"0008000004002040000200100000000042800584488000103081880008800000",
INIT_04 => X"00005842802AC210001000000800001000004080100040140080040800003100",
INIT_05 => X"0400000040000080410800010001002000000000004000002010000040002000",
INIT_06 => X"10100001221911E1911902000020200201A2D3E8000C2C84880010080800004C",
INIT_07 => X"C0002204000200000B080000010C040004A0400000C0000810000C5901036000",
INIT_08 => X"002A84300000014000C2008088090000002000000000030F8000001220000408",
INIT_09 => X"210000020000120082088801080020400000084010002880000C803400000008",
INIT_0A => X"020000040000480100D0010019019190200008B2022380800802010000000801",
INIT_0B => X"09000119064C810500D0A36851B428DA14368C801A1400000100500400000090",
INIT_0C => X"08100080000000A00000100080000000A00000000212000000000000B0001000",
INIT_0D => X"00100400000000A00000100400000000A0000540000000000000000000005100",
INIT_0E => X"00000000A8000900000040000000000000060000420000010000000000000120",
INIT_0F => X"4000040000102000000000020000000000000000240000800140000000000000",
INIT_10 => X"00001204FC000000000000000001280013A000400000000900E8000400000002",
INIT_11 => X"0000000001480004D5800004000000000000091D008000000000480740200000",
INIT_12 => X"0002000000000000000820080004DD000000000000000002A00011DC00001000",
INIT_13 => X"0322C01032301006022082000010032024200000048019500000000832901A80",
INIT_14 => X"4501000200089400007200D0020008000000144C4800000200BC228404020080",
INIT_15 => X"0010000104001000010440080000822900000000801010500A13404111008000",
INIT_16 => X"D1A0CA0000984D06403600086591900224002000400440104001040010000104",
INIT_17 => X"8DA368DA3685A1685A1685A1685A1685A1685A1685A1685A1685A1685A120D08",
INIT_18 => X"5A1685A1685A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA36",
INIT_19 => X"000000000000685A168DA368DA368DA368DA368DA368DA368DA368DA1685A168",
INIT_1A => X"6C20080AB9A28724904120E1999E91BCD151200802001038E2550A0010100000",
INIT_1B => X"68341A0D14514514514514514514514514514514514514534D34D34D34D344A1",
INIT_1C => X"268341A0D069349A0D069349A0D068341A4D268341A4D268341A0D068341A0D0",
INIT_1D => X"00000000000000000000000000000000000003FFFFFFFFFFFFFF8A6AC8341A4D",
INIT_1E => X"C2000557FEABEFA2D1400AA5D2AAAA00F7FFEAA10F7D17FFFFAAAE8000000000",
INIT_1F => X"03DFEFF7FFE8ABAF7802ABEFAAAE820000000021EFAA843DE00F7803FEBAFFFF",
INIT_20 => X"843DE00557BEAABAA2AEAABEFF78015555AA80174105555421EFF78028BEF5D0",
INIT_21 => X"504175FF0851401455555555EFA2FBC01FFF7AAAAB45557BC0155007FFDEBAAA",
INIT_22 => X"552A974AAA2843DEAA5D2A820BA000428AAAAA84154AAA2AA955FF00043DE005",
INIT_23 => X"AF7D1400BAAAAE821EFF7D17DEAA5D2AAAAAA5D557DE105D2EBDF55557FFDE00",
INIT_24 => X"BAFF803DF45FFD17DFFFFFD56AA00557FC201000517FFEFAAAEBDF45FFAEA8AB",
INIT_25 => X"FD7A2A48000000000000000000000000000000000000000000002ABFFA280154",
INIT_26 => X"AE38FF843DEBAEBFFC20285D75EFBC7A2DB400824120ADA38E3F1EFA28F7DF7D",
INIT_27 => X"421C7FF8028BEF41003FFD7F7F1EDA82F78E2DBD7A2A482038000A001C7A2803",
INIT_28 => X"1C716D1475FFEAAA28E3FE385D71E8AAAAAA0A8BC7EB8417555AA84104385D55",
INIT_29 => X"AA955C708003FE285D00155FF0055451555D5F575C7A2FBC51EFEBA0A8B6D557",
INIT_2A => X"12EBFF45497FFFE105D2E97482AA8038EAA412E850AA1C0428ABAB68E124BAA2",
INIT_2B => X"B6A0BFF55F7AEAAA82FFDF40092B6A4871EFFFD57FE825520ADA92495B7AE104",
INIT_2C => X"0000028BEFA28E124AAF7843AF7DEBDB78FFFE3DF6DA284175C001000557FFEF",
INIT_2D => X"AAA2D57FEAAF7FBFDF45AA800000000000000000000000000000000000000000",
INIT_2E => X"0BA082E82155AA802AAAAFF803DEBAAAFBC20BA55517DF55A2FBC201008003DE",
INIT_2F => X"5545A284000BA5D5340145F78028BFF08003DF45FFD57FE00FFAABFF45AA8002",
INIT_30 => X"D75FFA2842ABFF5555575FF55557FEAAA2AABFEAA5D5568ABAA2842AB55A2801",
INIT_31 => X"028ABAF7AA820BAAAAE9754500043DEBA5D04175EF0855575455D7BD5555A2FB",
INIT_32 => X"003DE00007FEAA10002ABFF450079FFE005D2A97400A2802AABA002A954AA5D0",
INIT_33 => X"0514200008517DFEFFF803FF45FFAAA8A00F7FBC2010FF80155EFF7D57DE005D",
INIT_34 => X"000000000000000000000028BFFA2AE820AAFF802ABEFAAFFEABEFAAFFFDEAA0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000200000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110204",
INIT_02 => X"0801080200100000046558040080000041000000002402400800000009008010",
INIT_03 => X"00020201040000D0842242024210810802006400088000003080054288C10000",
INIT_04 => X"0000400088020000003020002000001002A0E881108032100002000800203040",
INIT_05 => X"04092A081000411841480001000000201000012800400010001081C040402000",
INIT_06 => X"10100001220001E0001802002020240208000369001520080100100909000266",
INIT_07 => X"4000220440020000090C0810210A040004A0410000C0000810000C4901036008",
INIT_08 => X"0000802100100140004200808809000C002000000000010F8102041320000000",
INIT_09 => X"2000000000000200828888800808000410800840100220211850004442004048",
INIT_0A => X"240A80800442400004C0010000060210200008B2022304880800410000200801",
INIT_0B => X"0000010008008020020100008000400120800004004821202001A05A00040180",
INIT_0C => X"08101400000000A01004101400000000A0100000081300410402080080003000",
INIT_0D => X"04101080000000A01004101080000000A0100540000040000000000000405100",
INIT_0E => X"00000040A80009000180000000000000004608004200040800000000000001A0",
INIT_0F => X"4000282000102000000080008000000000000000240800800140000040000000",
INIT_10 => X"00001A00000002000000000020013000100010080000000D0000040040000003",
INIT_11 => X"0000000021500000800010400000000000400900000088000000680000009000",
INIT_12 => X"008000800000000000086010000080000100000000000082C000100000200800",
INIT_13 => X"040004924040008020000200101100004000000000C019500050000800000000",
INIT_14 => X"4541008240801000804000108280800001001051A12481041080801010000080",
INIT_15 => X"4800048004480044800044000240022100884000901210440003C141102B088A",
INIT_16 => X"00044280009048485D4020080000140004046240020044000480044800448000",
INIT_17 => X"080200802008020080200802008020080200802008020080200802048026E011",
INIT_18 => X"0000000000000000000000000002008020080200802008020080200802008020",
INIT_19 => X"0000000000000080200000000000000000000000000000000000000000000000",
INIT_1A => X"CA83332A34488A8A28A29E195281FC1A72E24C2BF5A4D9555204428290100000",
INIT_1B => X"94CA65328A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A354",
INIT_1C => X"994CA6532995CAE572B94CA6532994CA6572B95CAE532994CA6532994CA65329",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF838CF1CAE532",
INIT_1E => X"7FFFFAAAE801FF08557DF4555516AA00007BEABEFAAD1555FFF7840000000000",
INIT_1F => X"56AA0000043FFEFA2FFFDE1008556ABEFA2D1400AA5D2AAAA00F7FFEAA10F7D1",
INIT_20 => X"84020000000021EFAA843DE00F7803FEBAFFFFC2000557FC0010AAD57FF45A2D",
INIT_21 => X"7FFE8ABAF7802ABEFAAAEA8BFF5D0415400F7FBFDEAA007FEAB45AAAE800AAF7",
INIT_22 => X"5D0415555557BFDFEF00517DE00A28028B450855421EFF78028BEF5D003DFEFF",
INIT_23 => X"A5D7FFDEBAF7AEBDE00557BEAABAA2AEAABEFF78015555AA80174105555401FF",
INIT_24 => X"FFF7AAAAB45557BC0155007FFDEBAAA8417410AAFFD7555AAD56AB45A2AE800A",
INIT_25 => X"5C7E380000000000000000000000000000000000000000000000155EFA2FBC01",
INIT_26 => X"DA38E3F1EFA28F7DF7DFD7A2A4801EF085F7AF6D55556AA381C75EABEFBED157",
INIT_27 => X"C0010AADF7AF6DB6D56FA3814003AFFFA2F1F8E381C516FBC7A2DB400824120A",
INIT_28 => X"5E8B45BEA0850BAE38002038000A001C7A2803AE38FF843DEBAEBFFC20285D75",
INIT_29 => X"8028BEF41003FFD7F7F1EDA82F78E2DBD7A2A4ADBEF550412428F7F5FDE92087",
INIT_2A => X"A84104385D55401C75504125455575FAFD7145578E10AA802FB450851421C7FF",
INIT_2B => X"BED56FB45BEA082082557BF8EBAF7AABFE385D71E8AAAAAA0A8BC7EB8417555A",
INIT_2C => X"00000175C7A2FBC51EFEBA0A8B6D5571C716D1475FFEAAA28E10438AAF5D2545",
INIT_2D => X"BA5D5568BEFF7D157555AA800000000000000000000000000000000000000000",
INIT_2E => X"F55A2FBC201008003DEAAA2D57FEAAF7FBFDF45AA80021FF007BE8BFF5D516AA",
INIT_2F => X"DEBAAAFBC20BA555140010AAFFE8BFFFFD17DEBA5D002ABFFA2D16AAAA55517D",
INIT_30 => X"020BAFFD17DE10005568B55FF80154BAA280020BA082E82155AA802AAAAFF803",
INIT_31 => X"43FF55085140145F78028BFF08003DF45FFD57FE00FFAABFF45AA803FFEF5500",
INIT_32 => X"842AB55A28015545A284000BA5D53421455504021555D556AB555D5568A00AA8",
INIT_33 => X"2AA800AAAAD142155F7D57DF45FF8002010557FEAAAAF7AABFEAA5D5568ABAA2",
INIT_34 => X"000000000000000000000015555A2FBD75FFA2842ABFF5555575FF55557FEAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000023FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B83008481800E0000C26426040000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"00080D4912E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"000048048002400048150000000002504230C899109032100020160880223000",
INIT_05 => X"040B2A229100410041088011100022201200012840440000B01088C0005C2400",
INIT_06 => X"287E4003225021C5021880C02000A40249048363A5992808110010090908022A",
INIT_07 => X"4044222987020C80152D8910210A0400252B74200045C86810000C5B0503286A",
INIT_08 => X"26509804400501400242C0B0B83B0134702000000000191FA162841324832069",
INIT_09 => X"3002000220001240820F8B2A08000040409018401001200159D80D64AA004041",
INIT_0A => X"020808852000420718C00101B0070310200008B60A23A51B2802467327200801",
INIT_0B => X"080802500C08832582810240812040912094068010050402214850444091019B",
INIT_0C => X"761B011986695014A96E1A8119865A5018C5A0A00012004104020808B0003000",
INIT_0D => X"AE1A811986695014A96E1B0119865A5018C5AF0062C38A4DB680A0D8241501D5",
INIT_0E => X"802CAB184E8F4101621B1BAC845542056A289A1BB2078A922DA2A8B180A2600A",
INIT_0F => X"392000224ACDE215883078681B5C05AA429189B60AC43CEC7F0272C3841DB528",
INIT_10 => X"51BCA1C90006C0C2958502861120C003104289A668B8CAB270106338317A3D94",
INIT_11 => X"A64090B89E015AAA880E48382EB8804B020A06020C67061BC785938085134CD5",
INIT_12 => X"C6284B2D20410AB4503089C00A8280819A5539D503336D61056ABA006282806C",
INIT_13 => X"060040142020015001004A00080042004000E8089C9003066E03513E41470126",
INIT_14 => X"4536708201C000908020349320008000A1000C09A9348498B000000000000080",
INIT_15 => X"32A0C32A0C32A0832A0C19504195040040000000801010028001400010010CBA",
INIT_16 => X"8104400000904C0C0964200841010954000444D280140050C32A0832A0C32A08",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090246811",
INIT_18 => X"1004010040100401004010040102409024090240902409024090240902409024",
INIT_19 => X"0000000000004010040100401004010040100401004010040100401004010040",
INIT_1A => X"488292A831308E0000000A11100830181621409A14E871104201400284000000",
INIT_1B => X"0000000000000000000000000000000000000000000000020820820820820A05",
INIT_1C => X"0000000402000000000000000000010080000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8C0F00000000",
INIT_1E => X"555FFF784020AAF7D542155F7D1400AAF7FFFDE00F7842AA00002A8000000000",
INIT_1F => X"A800AA007FFDFFFA28428A000000001FF08557DF4555516AA00007BEABEFAAD1",
INIT_20 => X"FBEABEFA2D1400AA5D2AAAA00F7FFEAA10F7D17FFFFAAAEA8ABAFFD17FEBAFFA",
INIT_21 => X"0043FFEFA2FFFDE1008556AB45555568A10A2FFC00AAF78028AAAFF84020AAFF",
INIT_22 => X"FFD1555FF0804000AA000428A10AAAA801EFFFD140010AAD57FF45A2D56AA000",
INIT_23 => X"FA2FBFFF550000020000000021EFAA843DE00F7803FEBAFFFFC2000557FC0155",
INIT_24 => X"00F7FBFDEAA007FEAB45AAAE800AAF78428B45A28428A10087FD7400552EBDFE",
INIT_25 => X"A101C2A80000000000000000000000000000000000000000000028BFF5D04154",
INIT_26 => X"AA381C75EABEFBED1575C7E380000BAF7DB4016DE3DF450AAF7F1FDE38FF8A2D",
INIT_27 => X"AFABAFFDF7AE82F7AA870AA0071F8FFFBE842DA101C0E001EF085F7AF6D55556",
INIT_28 => X"42DAAAE38A02082E3FBEFBC7A2DB400824120ADA38E3F1EFA28F7DF7DFD7A2A4",
INIT_29 => X"DF7AF6DB6D56FA3814003AFFFA2F1F8E381C516DB455D5B68A28A2FFC20AAEB8",
INIT_2A => X"BFFC20285D75C2145F7DF525EF140A050AA1C0028A28AAA4801FFE3DF40010AA",
INIT_2B => X"007FD74284120BFFFFBEF1F8F7D080A02038000A001C7A2803AE38FF843DEBAE",
INIT_2C => X"000002DBEF550412428F7F5FDE920875E8B45BEA0850BAE3802DB6DAA8A28A00",
INIT_2D => X"AAF7D57DEAAF7AABDE10552E8000000000000000000000000000000000000000",
INIT_2E => X"1FF007BE8BFF5D516AABA5D5568BEFF7D157555AA80020BAFFFBC01EFA2FFD74",
INIT_2F => X"FEAAF7FBFDF45AA803FEBAFFFBEAA00F7AE974BA085568BEFF7803FE10552E82",
INIT_30 => X"EAAAAA2FFC00AAAA803FEAAA2AA82000A2FFFDF55A2FBC201008003DEAAA2D57",
INIT_31 => X"0001FFAAFFC0010AAFFE8BFFFFD17DEBA5D002ABFFA2D16AAAA55517DF55557F",
INIT_32 => X"802AAAAFF803DEBAAAFBC20BA555142155F7FFC01EF552E974BA550028ABAA28",
INIT_33 => X"2803FFFFA2AAAAA00007FD74BA08003DFFFFFD16ABFF082E820BA082E82155AA",
INIT_34 => X"00000000000000000000003FFEF5500020BAFFD17DE10005568B55FF80154BAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000200000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702684000000008000008820009280A553231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"421A0A0012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"02004000890200001837830011998C31C09060DC104000102002140900003548",
INIT_05 => X"0402002BC200009841090001200006200800000020480010A4100100001C2000",
INIT_06 => X"287FC003230001D0001806C0060CB0622000037085C820000000100C0C200008",
INIT_07 => X"CE64B663DFA314C803292140890C0601F472D1640051F80C10020C493F033432",
INIT_08 => X"67C081000111814004C20481A92940EA7A3020480000071F846890162E135038",
INIT_09 => X"240048108488024082488BAF08000020800629441004300421800F04F8000001",
INIT_0A => X"A0200E0BF40063FF9DC0010000180018200408B27E234913E900067F04D40C01",
INIT_0B => X"002002801000A04200000000000000000000029D204B7C0382FD0100F3F9F80F",
INIT_0C => X"7E0B348EDAC3900F6EFA0B158EDA93900F6EE230381208008001007A80001100",
INIT_0D => X"CA0B158EDAC3900F6EFA0B348EDA93900F6EE8421392C96B1237E0D8BD9628F9",
INIT_0E => X"412EDD2B47CFF812A383430C669E622DBC31D73F6006A5891533EF9500EAE64B",
INIT_0F => X"BA30E022DAD8C100CA39E8CEBE66C2B083798D341B10DE7E14400392C74CAEAD",
INIT_10 => X"71A9C5DD00B12728D5360234D62A49FAB442994B3238D4E2FB104636652E19B8",
INIT_11 => X"C800DA550C29F36A8A2554E48A6430469392526208C6CC95C33717D885329664",
INIT_12 => X"51B60585A5C28895962502E9F36A828C4999AF580395542D27CDBA0020F0FABA",
INIT_13 => X"0000001E404011F066000A000EE040000000873FB80B8A00EF03F56CC12B416A",
INIT_14 => X"4D667C06CC6816B300403C13E2000000460010400000010CE080801010000080",
INIT_15 => X"72F0C72F0872F0872F0C597863978421040800209010124ACA03414158228430",
INIT_16 => X"00104280A89A4D004000000800001D5E05182493C5BC5AF0872F0C72F0872F08",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000010000",
INIT_18 => X"8020080200802008020080200800000000000000000000000000000000000000",
INIT_19 => X"0000000000000080200802008020080200802008020080200802008020080200",
INIT_1A => X"E02000028DCA05A8A28A2048C1111026C152A2316246000CB054420210100000",
INIT_1B => X"C864321904104104104104104104104104104104104104124924924924924481",
INIT_1C => X"2C964B2592C964B2592C964B2592C964B2592C964B2592C964B2190C86432190",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800FFD64B259",
INIT_1E => X"2AA00002AAAA10FF8002155F7FFC2000080417555FFAA80155F7840000000000",
INIT_1F => X"FE8AAA080000155F7FFFDEAA0000020AAF7D542155F7D1400AAF7FFFDE00F784",
INIT_20 => X"2E801FF08557DF4555516AA00007BEABEFAAD1555FFF7842AB55080000145557",
INIT_21 => X"07FFDFFFA28428A00000028B4555043DFFFFFAE82000FF80020AAA2AAAABFF00",
INIT_22 => X"A284174AAFF8428AAAFF8415545AAFBD7545F7AAA8ABAFFD17FEBAFFAA800AA0",
INIT_23 => X"5F7FFFDEAA08556ABEFA2D1400AA5D2AAAA00F7FFEAA10F7D17FFFFAAAE80000",
INIT_24 => X"10A2FFC00AAF78028AAAFF84020AAFFFBC21550800000105D55400AA082A8215",
INIT_25 => X"145F7840000000000000000000000000000000000000000000002AB45555568A",
INIT_26 => X"50AAF7F1FDE38FF8A2DA101C2AAFA00EB8E0516DE3F5C000014041256DEBA487",
INIT_27 => X"2FB551C0E0516D417FEDA921C000017DEBF5FDE92080E000BAF7DB4016DE3DF4",
INIT_28 => X"0070BAAAAAADBD70820801EF085F7AF6D55556AA381C75EABEFBED1575C7E380",
INIT_29 => X"DF7AE82F7AA870AA0071F8FFFBE842DA101C0E2DB55410A3FFC7F7A087000FF8",
INIT_2A => X"7DF7DFD7A2A480000BE8A17482F78A28A92E3841556DA2FBD7545F7AAAFABAFF",
INIT_2B => X"41554508208208017DF7F5FDE9208556FBC7A2DB400824120ADA38E3F1EFA28F",
INIT_2C => X"000002DB455D5B68A28A2FFC20AAEB842DAAAE38A02082E3FBC217D1C0E05000",
INIT_2D => X"005504001FFAA8015545F7800000000000000000000000000000000000000000",
INIT_2E => X"0BAFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE10552EBDE00AAAE975FFAAD1420",
INIT_2F => X"8BEFF7D157555AA803DF45552E975EF007FFFE005504001FFAAD17DE00082E82",
INIT_30 => X"BFF55FF8017410FF84154BAAAAABFF450000021FF007BE8BFF5D516AABA5D556",
INIT_31 => X"BD5555F7AEBFEBAFFFBEAA00F7AE974BA085568BEFF7803FE10552EBDF45002E",
INIT_32 => X"003DEAAA2D57FEAAF7FBFDF45AA8002000FFAE95400F7AEA8A10A284175FFAAF",
INIT_33 => X"2FFC21EF552A954100851554000004021FFFFD17DE1008517DF55A2FBC201008",
INIT_34 => X"00000000000000000000003DF55557FEAAAAA2FFC00AAAA803FEAAA2AA82000A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00020201926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"00104884880A4400403000004800027102A0E88110D83210642EA809C0203040",
INIT_05 => X"04092A08138041184109C001380000201A008128044E00754010C9C192D82400",
INIT_06 => X"201800012372A1D72A180000204024024954A3670819290951001009092C0222",
INIT_07 => X"4000220B40020C80052C0A12292A040005715540015E006810001C4B01032C7E",
INIT_08 => X"9032881000140140024200808839005C002010800000155F8122851320016400",
INIT_09 => X"2C80080200801280825A988008000040008208401005B3071859006442004054",
INIT_0A => X"200810940400720005C0030192072310200028B6022346080802E001A5600801",
INIT_0B => X"206822F20CA8826AC2A14250A128509528954404144C200425010040000001B0",
INIT_0C => X"A41AA5B7344C10B383081BA4B7341C10B3831034081200000000000430003000",
INIT_0D => X"381BA4B7344C10B383081AA5B7341C10B383110218CB0E54C2EA404A4F03D404",
INIT_0E => X"A008E730A01AB113A5524E6ACA678001CE3E20A5B284ED1132909C72885A2B2C",
INIT_0F => X"6430202021252991C22C99731014AC3CC0C0B8182597A801610218CB0C3548B3",
INIT_10 => X"5194332B018A444AEA2701288A15A151EC5952E44128CA194517354C180A3C06",
INIT_11 => X"D50048A411C158BB0A7910142C771804C8A0ADA2E6A983014780CA28B2A5C882",
INIT_12 => X"F8BE8E3E1E0109472C3EB50158BB02D09852745F80112C428562EE0353635232",
INIT_13 => X"02414032646000826080C20001104240480068001C9B9150A0000297046E4023",
INIT_14 => X"4510008241C80290882400908000A000A1000809A93485D61000000000000080",
INIT_15 => X"00000000040000000000000020000000000000008010102A82014100101118BA",
INIT_16 => X"A10441010090480C096420184321040002844840000000004000000000400000",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094246A10",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"0000000000005094250942509425094250942509425094250942509425094250",
INIT_1A => X"BFBFBFBF7DDF3BAAAAAABEFDDFE7EFBEFFE7CFC3F7EFFF7DF7E24502A8000000",
INIT_1B => X"F5FAFD7EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAFFD",
INIT_1C => X"BF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EB",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800FFDFAFD7E",
INIT_1E => X"80155F7842AB55552E821FFFFD5555EF552ABDFEF007FE8A00AAFBC000000000",
INIT_1F => X"BD55EFAAD1554BA00556AA00AAD16AA10FF8002155F7FFC2000080417555FFAA",
INIT_20 => X"55420AAF7D542155F7D1400AAF7FFFDE00F7842AA00002A821EF5D7BC21FFFFF",
INIT_21 => X"80000155F7FFFDEAA00002AB45082A821EF5D557FF45A2AABFEBA082A975555D",
INIT_22 => X"A2FFE8BEF5D517FF455D554214500043DEBAAAFFEAB55080000145557FE8AAA0",
INIT_23 => X"0552EBFEAAAAD1401FF08557DF4555516AA00007BEABEFAAD1555FFF7842AABA",
INIT_24 => X"FFFFAE82000FF80020AAA2AAAABFF002E80000AAAABDF555D2E955EFA28428A1",
INIT_25 => X"A28AAF5C0000000000000000000000000000000000000000000028B4555043DF",
INIT_26 => X"000014041256DEBA487145F78428B6D4120851FFEBD5525C74124B8FC71C71EF",
INIT_27 => X"871C74975C01FFEBF5D25EFA2D555482085F6FA28AAD16FA00EB8E0516DE3F5C",
INIT_28 => X"0BFE921C2E9557D415B400BAF7DB4016DE3DF450AAF7F1FDE38FF8A2DA101C2A",
INIT_29 => X"0E0516D417FEDA921C000017DEBF5FDE92080E2AB7D1C24851FF495F7FF55A2A",
INIT_2A => X"ED1575C7E38028A82B6F1E8BFF495F78F7D49554214508003FEAABEFFEFB551C",
INIT_2B => X"5D20905C7AA842DA00492EBFEAABED1401EF085F7AF6D55556AA381C75EABEFB",
INIT_2C => X"000002DB55410A3FFC7F7A087000FF80070BAAAAAADBD7082087000AAA4BFF7D",
INIT_2D => X"4508042AB455D517DEBAA2D54000000000000000000000000000000000000000",
INIT_2E => X"E00AAAE975FFAAD1420005504001FFAA8015545F78028BFF0004175EFA2D5421",
INIT_2F => X"DEAAF7AABDE10552E975450051401EFA2D5421EFAAD557410007BFDEAAA2D57D",
INIT_30 => X"175FF087BFFF45AA843FE005D2A955FF087BC20BAFFFBC01EFA2FFD74AAF7D57",
INIT_31 => X"03FEBAFFFBFDF45552E975EF007FFFE005504001FFAAD17DE00082EA8BFF5504",
INIT_32 => X"516AABA5D5568BEFF7D157555AA8028A00FFD16ABFF087BEABEF005542155000",
INIT_33 => X"00017410AA803DFEF550402155A2843FE00082ABFEAAFFD5421FF007BE8BFF5D",
INIT_34 => X"00000000000000000000003DF45002EBFF55FF8017410FF84154BAAAAABFF450",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000033FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"0002074F200904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000480488024000403000000000001002A0E881108032100002000800203040",
INIT_05 => X"04092A081000411841080001000000201000012800400010001081C000402000",
INIT_06 => X"80500001221021C1021800002000240249048361001128081100100909000222",
INIT_07 => X"4000220050020480152D0A142D0A8400043B45400040006810000C5901033D78",
INIT_08 => X"0010880000100140024280808829029C002000000000053FA142051324902030",
INIT_09 => X"2000000000000200820888800800004000800840100020011858006442004040",
INIT_0A => X"200800840400400005C0010190070310200008B202236D080802400001600801",
INIT_0B => X"000000100C088020028102408120409120940404104C20002101004000000110",
INIT_0C => X"5210040000B0E0A0000210040000E0E0A0000190081200000000000000003000",
INIT_0D => X"0210008000B0E0A0000210008000E0E0A0000B02740421A0E5D1A02400205080",
INIT_0E => X"40110080A4006110510C14D18178E01200860008920106460D4501CB00011130",
INIT_0F => X"411420220080220C0093C38923240ABBC00905C33C6000400F02740412C0715C",
INIT_10 => X"8000120800658992F3C700C3018120000041DB011CC000090012565306500002",
INIT_11 => X"E240240A8340000200067EAA8CB65809240C09024A4AE0CA0000480083968239",
INIT_12 => X"7DB0D0200900422ACA4B28000002002B46867DBC002A830280000800F7B7A0B1",
INIT_13 => X"020040126060008020000200000042004005800004801150A00341244000845C",
INIT_14 => X"4500008240800000802000908000800001000009A92481041000000000000080",
INIT_15 => X"000040000000000000040000000000000000000080101000000141001001088A",
INIT_16 => X"810440000090480C096420084101040000044040000000004000040000000000",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090246810",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"0000000000004090240902409024090240902409024090240902409024090240",
INIT_1A => X"EFBBBBAABCDABF9E79E7BEF9CB91FE1EF7D3AEB9F3E6FF7DF650400280000000",
INIT_1B => X"FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7FC",
INIT_1C => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8FF000FE7F3F",
INIT_1E => X"E8A00AAFBE8BEFA2D568ABA00003DF555555574AAAAAEAAB45082E8000000000",
INIT_1F => X"02AABA555155400557BC2010557BEAB55552E821FFFFD5555EF552ABDFEF007F",
INIT_20 => X"002AA10FF8002155F7FFC2000080417555FFAA80155F78428AAA007FE8A10080",
INIT_21 => X"AD1554BA00556AA00AAD140145AA8028ABA002EBFFFF082EBDEBAA2D1420105D",
INIT_22 => X"A2AEA8A10080428A10FFAEBFFEF5D0428B45A2FFC21EF5D7BC21FFFFFBD55EFA",
INIT_23 => X"5F7FBC0010FFAA820AAF7D542155F7D1400AAF7FFFDE00F7842AA00002A80155",
INIT_24 => X"EF5D557FF45A2AABFEBA082A975555D55400BA005568A000000175FFF7D15554",
INIT_25 => X"B6D00248000000000000000000000000000000000000000000002AB45082A821",
INIT_26 => X"25C74124B8FC71C71EFA28AAF5E8BFFB6D56DA82000E38F6D4155504AAA2AEAA",
INIT_27 => X"28ABA147FEDA10080E2AAAA555552400417FC20005D75E8B6D4120851FFEBD55",
INIT_28 => X"4BAEAAB6DB4202849042FA00EB8E0516DE3F5C000014041256DEBA487145F784",
INIT_29 => X"75C01FFEBF5D25EFA2D555482085F6FA28AAD147155BE8028A82002EB8FC7002",
INIT_2A => X"F8A2DA101C2A80145B6AEA8A10080E2DA00F7A0BDFD7550428B55A2F1C71C749",
INIT_2B => X"0004175FFE3D15757DE3F5C0038FFAA800BAF7DB4016DE3DF450AAF7F1FDE38F",
INIT_2C => X"000002AB7D1C24851FF495F7FF55A2A0BFE921C2E9557D415B400AA00556DA00",
INIT_2D => X"EF0051400AAA2AAAABFF08000000000000000000000000000000000000000000",
INIT_2E => X"BFF0004175EFA2D54214508042AB455D517DEBAA2D568BEFFFD57FE10002AAAB",
INIT_2F => X"01FFAA8015545F78028AAA557FFFE00082EAAAAA5D5142000007BC20105D5568",
INIT_30 => X"28A00082EAAB45000028ABAFFFBC20AA08043DE00AAAE975FFAAD14200055040",
INIT_31 => X"02AB55AAD1575450051401EFA2D5421EFAAD557410007BFDEAAA2D557555FF80",
INIT_32 => X"FFD74AAF7D57DEAAF7AABDE10552E82155FFAAA8A10002ABFE00F7803FF555D0",
INIT_33 => X"87BC20AA00517DE000804175EFAAD1555EFA2D1420BAFFAE820BAFFFBC01EFA2",
INIT_34 => X"000000000000000000000028BFF5504175FF087BFFF45AA843FE005D2A955FF0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000100000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"000440009282000001100000000000100220C8811080321000000228002A3000",
INIT_05 => X"04092A0010004300418800510000A6201000012A64400000145080C000422000",
INIT_06 => X"00100001220001C00018821020402402080003772019200001001009090002AA",
INIT_07 => X"4000220000021840010C8912250A0400042044400040006810000C4901032B18",
INIT_08 => X"0022810000058140024280A0A8190004002030C00000016F8122041320000000",
INIT_09 => X"20000000000002C0820888008800000000800840100020011850004402004040",
INIT_0A => X"00080094000062000180010180060210200008B2022304080800400003E00801",
INIT_0B => X"0000000008008020020000000000000100800000000000002500004000000130",
INIT_0C => X"0010108000000000000010108000000000000230001200000000000420003000",
INIT_0D => X"0010140000000000000010140000000000000100000040000000000000000000",
INIT_0E => X"0000000000000100008040000000000000000000020000090000000000000000",
INIT_0F => X"0030002000406000000000068409014000000000000000000100000040000000",
INIT_10 => X"0000000800000201000800000000000000400048000000000010000440000000",
INIT_11 => X"00A0000000000002000000441108800000000002008008000000000080201000",
INIT_12 => X"0242038B82800000000000000002000001000000000000000000080000001844",
INIT_13 => X"000000100000000005C04A000000400000000000000001062000000400000000",
INIT_14 => X"4500008200800000800000100000800001000001A12480001000000000000080",
INIT_15 => X"000000000000000000040000200002000000000080101000004140001001088A",
INIT_16 => X"0004400000904808094020080000000000044040000000004000040000400004",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000046000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000400280000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000000000",
INIT_1E => X"AAB45082EBFE000004020AA552E80000F7FBC214555003DE10A2FBC000000000",
INIT_1F => X"BE8A10F7802AA0055003FE10007BE8BEFA2D568ABA00003DF555555574AAAAAE",
INIT_20 => X"AEAAB55552E821FFFFD5555EF552ABDFEF007FE8A00AAFBFDEBA555568BEFA2F",
INIT_21 => X"55155400557BC2010557BFFFEFA2FFC20005D2A955EFF78428BEFAAD17DF55AA",
INIT_22 => X"5D2AA8B45AAD57FF55A2FBC21FFA28415400FF8028AAA007FE8A1008002AABA5",
INIT_23 => X"A002E9740055516AA10FF8002155F7FFC2000080417555FFAA80155F7843DF45",
INIT_24 => X"BA002EBFFFF082EBDEBAA2D1420105D003FFFF08514200055002AA00AA802AAB",
INIT_25 => X"E28B6FFC0000000000000000000000000000000000000000000000145AA8028A",
INIT_26 => X"8F6D4155504AAA2AEAAB6D0024B8E381C0A00092412A87010E3F5C0145410E3D",
INIT_27 => X"F8EAA495F68BFFA2F1EFA38E38428A005D0038E28147FE8BFFB6D56DA82000E3",
INIT_28 => X"428BEFB6DB7DF45AAAEA8B6D4120851FFEBD5525C74124B8FC71C71EFA28AAF5",
INIT_29 => X"7FEDA10080E2AAAA555552400417FC20005D75F8FFFBEF5C0000492A955FFF78",
INIT_2A => X"BA487145F7843FF7D4120A8B6DAAD17FF55B6F5C21EFAA8E10400E38E28ABA14",
INIT_2B => X"41002FA38A2842AA82142095428415F6FA00EB8E0516DE3F5C000014041256DE",
INIT_2C => X"0000007155BE8028A82002EB8FC70024BAEAAB6DB4202849043FFC7005F45010",
INIT_2D => X"00A2D542155002ABDEBAF7FBC000000000000000000000000000000000000000",
INIT_2E => X"BEFFFD57FE10002AAABEF0051400AAA2AAAABFF08002AAAA5D2A82000082E954",
INIT_2F => X"AB455D517DEBAA2D56AABA087BEABEFAAD57DEAAA2802AA105D002AABA5D7BE8",
INIT_30 => X"42010082A955EFFF8428BFFFFFBFDF55A2AEA8BFF0004175EFA2D54214508042",
INIT_31 => X"A82000AAAAA8AAA557FFFE00082EAAAAA5D5142000007BC20105D556ABFFF7D1",
INIT_32 => X"D1420005504001FFAA8015545F7803FFEF08002ABEFA2D57DF45F7D1401FFA2A",
INIT_33 => X"8043FF55087BD740000043DEAAA2842AA005D00154AA007BFDE00AAAE975FFAA",
INIT_34 => X"000000000000000000000017555FF8028A00082EAAB45000028ABAFFFBC20AA0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000300000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"0202115002BB10080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"2FE962000017102918900948514522CE09200C0D590569398ADBF8CC1E50E480",
INIT_05 => X"5E6023002834854AE41C1E8782F508F2A15B71D412E0AFD9C2990DA56FF0B55A",
INIT_06 => X"B9B9E55402000340003200220A86012D0000000480D0400001555960540180A0",
INIT_07 => X"40D890101DBD400901442800817C2901F400868554DE240000A80090CE82A803",
INIT_08 => X"0122004000005665510320C9C90510025A8A00000A0A048F550A440E0001380C",
INIT_09 => X"2060410280081116C8204D016CB2CB290008008279580411289000000118A905",
INIT_0A => X"00008176802203180025699200140001A15000017F0051D0F837324E002A8A56",
INIT_0B => X"4485D000000124002400000000000001004010A8812831605DA0000A054052E4",
INIT_0C => X"B5320018CAC99BA0A3B9320018CAAAADA0C343F1AC1B01040A00202489551455",
INIT_0D => X"59320018CAC99BA0ACB9320018CAAAADA0CC421CA003B694B68018FAAA708E2C",
INIT_0E => X"B2449A3FF2FA04E5E09B128834ADB1443A1891E4A928C29020E6A8524CE7A3EE",
INIT_0F => X"2375B801324301AB0067622E5E5404B2A5A40B1E6644AF0F021EA003AC24352A",
INIT_10 => X"0A8C241815FEB6A9158863F638FB60ED838E890B703C6260D8E3A21275714C90",
INIT_11 => X"15F11133D171727A2550EE2F1BA0064F70DBDB1C74424E91E1C194C71D1216F5",
INIT_12 => X"432A2B2D001F803471A9A960E57245FDF9D364DBD9435A6D45C9E81BED555E4C",
INIT_13 => X"C00006B0800000038814B72AB01508150013F162119014204373517700ACCC59",
INIT_14 => X"300208092B940192D1000000000000A8A5AA80018120E00066000000000012CA",
INIT_15 => X"1000110001100011000108000880008000520228080108039501200848002912",
INIT_16 => X"081500008A422150884081AC9000010003561180063DB4F61100011000110001",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000012000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"BCBF0F2C688A8D3CF3CF0A7A898D21B4C9838D3030EF5168A360400000000000",
INIT_1B => X"E9F47A7D345345345345345345345345345345345345345145145145145147A5",
INIT_1C => X"3E9F4FA3D1E8F47A3D1E8F47A3D1E9F4FA7D3E9F4FA7D3E9F4FA7D1E9F47A7D1",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800001F4FA7D",
INIT_1E => X"3DE10A2FBC21FFFFFBFDF45A2D56AB45FFFFD54BAFF80001FF002A8000000000",
INIT_1F => X"FFFE005D7BC0010002E954AA087FFFE000004020AA552E80000F7FBC21455500",
INIT_20 => X"FFE8BEFA2D568ABA00003DF555555574AAAAAEAAB45082E974BA5D7BFDF55A2F",
INIT_21 => X"7802AA0055003FE10007BC0000082A97400550017410FFD1555550000020BAAA",
INIT_22 => X"AAFBD74105504021FF5D2EAAABAFFFBD55FF002ABDEBA555568BEFA2FBE8A10F",
INIT_23 => X"0007FC00AA087FEAB55552E821FFFFD5555EF552ABDFEF007FE8A00AAFBD55EF",
INIT_24 => X"005D2A955EFF78428BEFAAD17DF55AAAE820AA5D517DF45AAFFFFEAAFFAABFE1",
INIT_25 => X"1FF08248000000000000000000000000000000000000000000003FFEFA2FFC20",
INIT_26 => X"7010E3F5C0145410E3DE28B6FFC21C7E3F1F8F55AADB6FB6DFFFBD54AAE38E02",
INIT_27 => X"92482497BFDF45AAFFF8E385D7BC5000002E904BA1C7FF8E381C0A00092412A8",
INIT_28 => X"B555450804070BABEF5E8BFFB6D56DA82000E38F6D4155504AAA2AEAAB6D0024",
INIT_29 => X"5F68BFFA2F1EFA38E38428A005D0038E28147FC2010142E90428490015400FFD",
INIT_2A => X"C71EFA28AAF5D25D7B6F1D54384904021FF5D2AADAAAFFF1D55FF002EB8EAA49",
INIT_2B => X"A2F1FDEAAEBAABDE001471C20921475E8B6D4120851FFEBD5525C74124B8FC71",
INIT_2C => X"0000038FFFBEF5C0000492A955FFF78428BEFB6DB7DF45AAAE820925D5B7DF45",
INIT_2D => X"EFF7FFD54AAAAAA801EF00000000000000000000000000000000000000000000",
INIT_2E => X"AAA5D2A82000082E95400A2D542155002ABDEBAF7FBC2145AAD568B45AAFBFFF",
INIT_2F => X"00AAA2AAAABFF080000000087BFDF55A2FFE8AAA557FD7410082A800AA557BEA",
INIT_30 => X"800BA080417400F7FBD75450800174AAFFD168BEFFFD57FE10002AAABEF00514",
INIT_31 => X"1575EF082EAAABA087BEABEFAAD57DEAAA2802AA105D002AABA5D7BC20005D2E",
INIT_32 => X"D54214508042AB455D517DEBAA2D540155F7D1554AA0800001EF5D2ABDEBAF7D",
INIT_33 => X"2AE82010557FFDF55A2D57FEAAAAAEBFE10555140000555568BFF0004175EFA2",
INIT_34 => X"00000000000000000000002ABFFF7D142010082A955EFFF8428BFFFFFBFDF55A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000100000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"5295B6957FCBE0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"6DE90201BF90102103AF158E805428249851BFB2C106592088DBF8400A5055C2",
INIT_05 => X"3824BD7F80148D9E07100A8201ED01C1A19B68F40A807ED9C18114956FF081DB",
INIT_06 => X"6A8F033DD800000000050716BE9F57F8AC000807DFD9B00000CF20E5E1818B1B",
INIT_07 => X"86481240FE05A109228E2C0891D772A6F40045B8CF30E085DD2ED57D4EED08CA",
INIT_08 => X"DF23800005981C0338190549C904182B6113870022000488C08B46268A001508",
INIT_09 => X"823DF78CDB6CA60E0E28EFFE2061872F80C1684A80C8604085F0074D3B72637F",
INIT_0A => X"BD2FAD7FE653C3BA1FF33E0E001E000B3A5DAADAFDDA5DA79350CFB8013E7437",
INIT_0B => X"C5C3D00018006C681700000000000000020012E9E10A31EB5FF9296A67F5B4FF",
INIT_0C => X"542A6FEEB2533EA160782A6FEEB2333EA16031F2BD47BDA2CA5D8164FCCFE833",
INIT_0D => X"F82A6FEEB2533EA160782A6FEEB2333EA160391BEFF2C32FB695F919110D5ECE",
INIT_0E => X"5A86840354D1706FFFA3EF6E24B6D18C0D06638A207CFDE1F7DDAD76D5282400",
INIT_0F => X"4D77FAAB77CE3AF3EE78F58DB737E6E43E59AFE4A59B57679D19EFF2C7573FAD",
INIT_10 => X"72CA52606DFED6CA55334C04C04FF7D7A0ABD6DAAAB96529382B74E4E1FE4ACA",
INIT_11 => X"AA1A184045D5D7A870D2F5A5D7522D1281017F056E9C9C3FC95949C157ADB555",
INIT_12 => X"A58949D5B5C85F97871876F7D7E859FDEB974F486905001FDF5FA0D719F9956E",
INIT_13 => X"70021EE341036BF368128419FB5560158015177F916A039EF41FDB34A91F432E",
INIT_14 => X"1D0A7CC9AE7A08BFF0001D35682AC0CE8FCCC200A59BDD2FFE3F3EC7C7DEF206",
INIT_15 => X"BCF4FBCF4FBCF4FBCF4FBE7A7DE7A7800617112E46F05D02DD814102F800633F",
INIT_16 => X"00179C16DECF67F08BC02F9086000D9E8A3F06ABD73DBCF4FBCF4FBCF4FBCF4F",
INIT_17 => X"000000000000000000000000000000000000000000000000000000000005F080",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"930D0D1B9000303AEBAE88BE013DB9880A5D25C0408006114F981800C0000000",
INIT_1B => X"351A8D069A6BAE9A69A6BAE9A6BAE9A69A6BAE9A6BAE9A69A69A69A69A69A918",
INIT_1C => X"A351A8D46A351A8D46A351A8D46A341A0D068341A0D068341A0D068351A8D068",
INIT_1D => X"00000000000000000000000000000000000003FFFFFFFFFFFFFF8000011A8D46",
INIT_1E => X"001FF002A821FFFFFFFFFFFFFFBFDFEFAAD142010007BEAB55FFAA8000000000",
INIT_1F => X"A975EFA2D140145007BC21FF5D2A821FFFFFBFDF45A2D56AB45FFFFD54BAFF80",
INIT_20 => X"7BFFE000004020AA552E80000F7FBC214555003DE10A2FBEAB45A28000010082",
INIT_21 => X"D7BC0010002E954AA087FD7400082E954AA0800154AA0855575FFAAD57FE005D",
INIT_22 => X"F7D16AB45FFFFEABEF007BD74005555555EFF7AE974BA5D7BFDF55A2FFFFE005",
INIT_23 => X"5555568B45552EA8BEFA2D568ABA00003DF555555574AAAAAEAAB45082EBFFFF",
INIT_24 => X"00550017410FFD1555550000020BAAAFFC0145AA84154BA082E801FFAAFBC015",
INIT_25 => X"B7DEBA480000000000000000000000000000000000000000000000000082A974",
INIT_26 => X"FB6DFFFBD54AAE38E021FF0824851FFFFFFFFFEFF7F1FAFD7A2D5400001C7BED",
INIT_27 => X"EFB45AA8E070281C20925FFBEDB451451C7BC01EF4124821C7E3F1F8F55AADB6",
INIT_28 => X"5505EFBEDB7AE385D7FF8E381C0A00092412A87010E3F5C0145410E3DE28B6FF",
INIT_29 => X"7BFDF45AAFFF8E385D7BC5000002E904BA1C7FD54280024924AA1404174AA005",
INIT_2A => X"2AEAAB6D0024BFFD7FFDB6AB7DFFF5EDBC71C7BD54005D5B575EFEBAE9248249",
INIT_2B => X"1C20801FFB6F5C0145555B68B7D4124A8BFFB6D56DA82000E38F6D4155504AAA",
INIT_2C => X"0000002010142E90428490015400FFDB555450804070BABEF5C516DAA8A12492",
INIT_2D => X"45AAD5400005D7BFFFEFAA800000000000000000000000000000000000000000",
INIT_2E => X"145AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF0000155FFF7FBFDFEFFFD568B",
INIT_2F => X"2155002ABDEBAF7FBFDF55A2AA974AA5D04001EFFFFFD5545557BC21FF080002",
INIT_30 => X"000AA5500174AA0855421FFFFFBEAAAA5D7BEAAAA5D2A82000082E95400A2D54",
INIT_31 => X"BD75FFAAAA80000087BFDF55A2FFE8AAA557FD7410082A800AA557BD74BA0004",
INIT_32 => X"2AAABEF0051400AAA2AAAABFF08003FF55F7FFEABFFF7D57FF455D7FD54105D7",
INIT_33 => X"FD1555FFA2AA800105504001EFFFD140145557BE8BEF000028BEFFFD57FE1000",
INIT_34 => X"0000000000000000000000020005D2E800BA080417400F7FBD75450800174AAF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000033FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"080BA868803F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"42016B0C401F58495C900A4859552A611D9A640F5903B2388004004C08A06008",
INIT_05 => X"16226B107811422A641C08038040007060E0032801E0202000991B708280B501",
INIT_06 => X"B3B8E0FC86142B4142B0000000011114D305824024090A1A143F182000000000",
INIT_07 => X"802102401015610A02C4005000EA019D002482043FCF1C8090C02800C0120886",
INIT_08 => X"20D40A5004003260F9810541494D403D9B98810A0002C601000054B94A006880",
INIT_09 => X"6070000504102805C820C8016C30C250080C0182183804012A0A102200110180",
INIT_0A => X"E000108010230445A800FD865421432121804021C20452880C2D100000022E0C",
INIT_0B => X"C2060014250B9080008306C18360C1B0609C05013065CC042004040808084001",
INIT_0C => X"8582081483ACC15F9C3982081483CCC15F9CBA45505640000A402019003F140F",
INIT_0D => X"F982081483ACC15F9F3982081483CCC15F9FB1962FCB69E08AAAEAEBCDDF7C72",
INIT_0E => X"E3F8E7F5E3AC3620805298B15A3FEBF1CFFF7670ACC3811A28AB57523CDFEBFB",
INIT_0F => X"DC4041D4CF03138DD865103EFEEAC9002BF05800D875E63CC9962FCB52CAA02F",
INIT_10 => X"8DB7BFE25208E8F46A228BF8A757F1B72A8A800B7546DB9F1CA320037F01BD67",
INIT_11 => X"9509EAAE7FD3B749471C48F8A45981CCFAFDBF9464006FD037AEFAE5150016EA",
INIT_12 => X"8802A3AF8E8FB0440CE78773B709641256EC844B8AF92FD7CEDC24A9E181A8A2",
INIT_13 => X"C284601C2864000080113307E4800297D086E00036D2440E0880AAD62BEFF577",
INIT_14 => X"A88DCC2211E44174112840880000060D7030C30B885200D274004008080003C1",
INIT_15 => X"0308003080030800308001840018400400602A01880980037109700C04C44C92",
INIT_16 => X"8340000020301805002D008CD943626111C0D95C20C2030A0030800308003080",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B0680834",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"00000000000041B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1",
INIT_1A => X"60B22A145DF60B8208209679D701DC2E784601F95163897DF160000000000000",
INIT_1B => X"944A2512AAA8A28A28A2AAAAAA8A28A28A2AAAAAA8A28A28A28A28A28A28A244",
INIT_1C => X"8944A25128944A25128944A25128944A25128944A25128944A25128954AA552A",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8000004A2512",
INIT_1E => X"EAB55FFAA821FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E820BA55000000000000",
INIT_1F => X"16AB55A2D542000A2D5400BA0800021FFFFFFFFFFFFFFBFDFEFAAD142010007B",
INIT_20 => X"80021FFFFFBFDF45A2D56AB45FFFFD54BAFF80001FF002A821FFFFFFFFFEFF7D",
INIT_21 => X"2D140145007BC21FF5D2AAABFFF7D168B45AAD57DFFFFFFFC0010F7842AA10F7",
INIT_22 => X"000002010552E95410AAFBD75FF5D7FEAB5500516AB45A28000010082A975EFA",
INIT_23 => X"5A284155FF5D517FE000004020AA552E80000F7FBC214555003DE10A2FBEAA00",
INIT_24 => X"AA0800154AA0855575FFAAD57FE005D7BD74000804174AA5D00020BA55554214",
INIT_25 => X"0AA490A00000000000000000000000000000000000000000000017400082E954",
INIT_26 => X"AFD7A2D5400001C7BEDB7DEBA4871FFFFFFFFFFFFFFFFDFEFF7FFD74AA552A82",
INIT_27 => X"821FFF7F1F8FC7EBD568B7DB6DF47000AADF400AA080A051FFFFFFFFFEFF7F1F",
INIT_28 => X"1C2000F78A2DA38E38A021C7E3F1F8F55AADB6FB6DFFFBD54AAE38E021FF0824",
INIT_29 => X"8E070281C20925FFBEDB451451C7BC01EF4124ADBC7E3D56AB7DB6DF78FD7EBF",
INIT_2A => X"10E3DE28B6FFE8A101C0E05010412495428AAF1D25EF497FEAB7D145B6FB45AA",
INIT_2B => X"5D0A000BA555F47145BE8A105EF555178E381C0A00092412A87010E3F5C01454",
INIT_2C => X"00000154280024924AA1404174AA0055505EFBEDB7AE385D7FD7438140012482",
INIT_2D => X"EFFFFBD54BA5D2A820AA082A8000000000000000000000000000000000000000",
INIT_2E => X"5FFF7FBFDFEFFFD568B45AAD5400005D7BFFFEFAA80155FFFFFFFFFFFF7FBFDF",
INIT_2F => X"54AAAAAA801EF0000021EFF7D16AB55A2D56ABEFF7FBD5410AAFBC00AA002A95",
INIT_30 => X"68BFFF7FFEAB45AAD140010F7AABFEBAAAAA82145AAD568B45AAFBFFFEFF7FFD",
INIT_31 => X"BE8BFF557BFDF55A2AA974AA5D04001EFFFFFD5545557BC21FF08003FF55AAD1",
INIT_32 => X"2E95400A2D542155002ABDEBAF7FBE8A00552E954100000154AAA2D1421FF007",
INIT_33 => X"D7BD74BA5D0002010552E820AA5D7BD7545F7AA801EF55516AAAA5D2A8200008",
INIT_34 => X"0000000000000000000000174BA0004000AA5500174AA0855421FFFFFBEAAAA5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000100000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000010228001000000000000000000024001620280000000000354200004008",
INIT_04 => X"00016200001310090090004840004152C7208802590000388000004C08006000",
INIT_05 => X"1621008008100002641C0803804000702000000000E02000009900000000B100",
INIT_06 => X"0210200C00000000000000000000000080000000000000000003182000000000",
INIT_07 => X"C00D267001B880080700285020020AC98820022802400480405008901100A001",
INIT_08 => X"000000000000106009872048400C4000010D000008000204150A00815A010084",
INIT_09 => X"0000000000000004C80000002C30C200000000021808005800000000000E0E00",
INIT_0A => X"0000000000000000080025860000000080A00020602040800000000000022A04",
INIT_0B => X"C002000000000000000000000000000000000000000000000000000084000760",
INIT_0C => X"385598035D0008A003B05598035D0008A0034078104B41A41000000000031400",
INIT_0D => X"505598035D0008A000B05598035D0008A0004263C0343EDD414004042228DC0D",
INIT_0E => X"0401180DE053A98F6ECC739D8140040231068187C39F5A4F985C008902041124",
INIT_0F => X"227848D4303807FC8CC5508AEAED1BFBD406451B02000E033263C0343CB74050",
INIT_10 => X"00000018A700FCF980CC300318A2420851546B2400000040D8549B5800000010",
INIT_11 => X"40E40511802208D6B30C48F8A8A452210402120A936B0000000004C2A8D64800",
INIT_12 => X"0006362A2B6424287B08286208D6B1427ED430B41402D025082359700181C211",
INIT_13 => X"40000000000000000010030060009C000018440021011821B35254E99AF9E941",
INIT_14 => X"002000044000000000000000000002F0001F00002024B20002000000000002C0",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000040",
INIT_16 => X"00000000000000000000008C8000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"441189B9045D82A69A69803F47E18E0218CC0140400200441920000000000000",
INIT_1B => X"4C261309861861861A69861861861861A69861861861861861861861861861A1",
INIT_1C => X"84C26130984C26130984C26130984C26130984C26130984C261349A4C2613098",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000261309",
INIT_1E => X"820BA55003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A800105D2E8000000000",
INIT_1F => X"FFDFEFF7FFD54BA5D2EA8BFFFF84021FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E",
INIT_20 => X"AE821FFFFFFFFFFFFFFBFDFEFAAD142010007BEAB55FFAABDFFFFFFFFFFFFFFF",
INIT_21 => X"2D542000A2D5400BA08003DFFFFFFFFFFFFF7FBE8B55A2D540010007BEAABAA2",
INIT_22 => X"FFFFFDFEFA2D56AB45AAFBD74AAFFD5420100804021FFFFFFFFFEFF7D16AB55A",
INIT_23 => X"AFF802ABFFFFAE821FFFFFBFDF45A2D56AB45FFFFD54BAFF80001FF002ABDFFF",
INIT_24 => X"45AAD57DFFFFFFFC0010F7842AA10F780155FFF7FBE8B45AAD568BFFF7FBD74B",
INIT_25 => X"000412A8000000000000000000000000000000000000000000002ABFFF7D168B",
INIT_26 => X"DFEFF7FFD74AA552A820AA490A38FFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2A80",
INIT_27 => X"BAFFFFFFFFFFFFF7FBFDFD7EBF1D24AA5D2AADBD7E384071FFFFFFFFFFFFFFFF",
INIT_28 => X"140000007FEFA92A2AA851FFFFFFFFFEFF7F1FAFD7A2D5400001C7BEDB7DEBA4",
INIT_29 => X"F1F8FC7EBD568B7DB6DF47000AADF400AA080A3FFFFFFFBFDFC7E3F5EAB45AAD",
INIT_2A => X"38E021FF0824BDFEFE3F1F8FD7AAD16DB7DBEFBD74AAE3DF400000004021FFF7",
INIT_2B => X"B6DB6FBD7E3F5D04AAFF8A2DBD7E3A0821C7E3F1F8F55AADB6FB6DFFFBD54AAE",
INIT_2C => X"000002DBC7E3D56AB7DB6DF78FD7EBF1C2000F78A2DA38E38A125C7E3F1EAB55",
INIT_2D => X"FFF7FBD54BA552A80010002A8000000000000000000000000000000000000000",
INIT_2E => X"5FFFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA082AA8BFFFFFFFFFFFFFFFFFF",
INIT_2F => X"00005D7BFFFEFAA8028BFFFFFFFDFEFF7FFFFF55A2D5400AA552ABDF55A28015",
INIT_30 => X"FDF55AAD16AB55AAD140010007BFFE10AAAA955FFF7FBFDFEFFFD568B45AAD54",
INIT_31 => X"BC20100800021EFF7D16AB55A2D56ABEFF7FBD5410AAFBC00AA002ABDFEFF7FB",
INIT_32 => X"FBFFFEFF7FFD54AAAAAA801EF00003FFEFA2D56AB45A2D57DFFFFFFFD54AAA2F",
INIT_33 => X"AAA82155AAD568B55FFFFFDF55A2D1400AAF7AABFF45AA8002145AAD568B45AA",
INIT_34 => X"00000000000000000000003FF55AAD168BFFF7FFEAB45AAD140010F7AABFEBAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000200000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"0001E6000053300B00D0005800000000000000407B0004BB830004DC3D01E000",
INIT_05 => X"FEE0000008720043EC3C3D0F87FA19F7E0201C409BE1F10623BB000A100CF300",
INIT_06 => X"06102FFC8E0007C00078008000171175A200096404D9404003FFDBE4744200AA",
INIT_07 => X"482491301000010001DC00000000000000004203FE4005800000008030002000",
INIT_08 => X"20E2008000027FEFF946058180010429000001080AAA010F8000000000000000",
INIT_09 => X"400000120000913FD80000003DF7DE0080010047FBF8000000000800C5408000",
INIT_0A => X"0080000010000400080FFDBE000000400000010000010050600220461003EAFE",
INIT_0B => X"C00600000000801020000000000000010240001721214E000004000000080000",
INIT_0C => X"08020000200000000F30020000200000000F3008001E00000000001803FF14FF",
INIT_0D => X"F0020000200000000F30020000200000000F3040200000020000000026A70C00",
INIT_0E => X"000019B140000800800000020000000030B86000400080000200000000004A58",
INIT_0F => X"AC08000000508001030A0A4001000000000002183E61E6000040200001000000",
INIT_10 => X"0000A56000090100000000001F86C00010080000000000525801000000000014",
INIT_11 => X"0000001716800000803102020000000002BC360020000000000292C010000000",
INIT_12 => X"DF70C08040100000706707600000801000000000000057450000100106060000",
INIT_13 => X"C011001C81080001101F977FE00800000000000040040040002000080506049C",
INIT_14 => X"0000000000000000020020029000000000000000020000000000000000000ADF",
INIT_15 => X"0000000000000000000000000000000000000000000002000200000000000000",
INIT_16 => X"0801810100000000000093ED8000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000401008080",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"930424038000343CF3CF349600704000201120A983400E0104D2040020000000",
INIT_1B => X"190C86432CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB0C30C30C30C30C818",
INIT_1C => X"2190C86432190C86432190C86432190C86432190C86432190C86432190C86432",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8000010C8643",
INIT_1E => X"800105D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8201008040000000000",
INIT_1F => X"FFFFFFFFFBD54BA552A8001000003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A",
INIT_20 => X"2E821FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E820BA5500001FFFFFFFFFFFFFF",
INIT_21 => X"7FFD54BA5D2EA8BFFFF843FFFFFFFFFFFFFFFFFFFFEFF7FFD74BA552E801FF00",
INIT_22 => X"FFFFFFFFFFFFBFDFEFFFD542000082EAAB55AAAABDFFFFFFFFFFFFFFFFFDFEFF",
INIT_23 => X"0087BE8B55F784021FFFFFFFFFFFFFFBFDFEFAAD142010007BEAB55FFAA801FF",
INIT_24 => X"FFF7FBE8B55A2D540010007BEAABAA2AE975FFFFFFFFFFFF7FBFDF55AAD14000",
INIT_25 => X"00014000000000000000000000000000000000000000000000003DFFFFFFFFFF",
INIT_26 => X"FFFFFFFBD54AA5D2A80000412ABFFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A82",
INIT_27 => X"021FFFFFFFFFFFFFFFFFFEFF7FBD74BA5D2A800281C0038FFFFFFFFFFFFFFFFF",
INIT_28 => X"FD54BA5D2A801C7142E871FFFFFFFFFFFFFFFFDFEFF7FFD74AA552A820AA490A",
INIT_29 => X"FFFFFFFF7FBFDFD7EBF1D24AA5D2AADBD7E38438FFFFFFFFFFFFFFFBFDFEFFFF",
INIT_2A => X"C7BEDB7DEBA4871FFFFFFFFFEFF7FBF8FD7E3D140010142AAFB7DBEAEBAFFFFF",
INIT_2B => X"E3F1FAF45A2D142010087FEDB55F78A051FFFFFFFFFEFF7F1FAFD7A2D5400001",
INIT_2C => X"000003FFFFFFFBFDFC7E3F5EAB45AAD140000007FEFA92A2AA925FFFFFFFDFEF",
INIT_2D => X"FFFFFFD74AA552A820005D040000000000000000000000000000000000000000",
INIT_2E => X"BFFFFFFFFFFFFFFFFFFFFF7FBD54BA552A80010002ABFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"54BA5D2A820AA082A821FFFFFFFFFFFFFFBFDFEFF7FFD74AA5D2A800BA550428",
INIT_30 => X"FFFEFF7FBFFFFFF7FBD74BA552A80145552E955FFFFFFFFFFFF7FBFDFEFFFFBD",
INIT_31 => X"ABFFFFFFAEA8BFFFFFFFDFEFF7FFFFF55A2D5400AA552ABDF55A2802ABFFFFFF",
INIT_32 => X"D568B45AAD5400005D7BFFFEFAA80175FFFFFBFDFEFF7FFEAB45AAD1420105D2",
INIT_33 => X"AAA821EFF7FBFDFFFAAD168B55A2D542010007BFDF55F7AE955FFF7FBFDFEFFF",
INIT_34 => X"00000000000000000000003DFEFF7FBFDF55AAD16AB55AAD140010007BFFE10A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"1094EC681244819000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"0001E6000053300F01D4587800446194F49020107F0012BBC00202DC3823EA82",
INIT_05 => X"FFF201B228704123FC3C381F87C03DFFF012412A9FE1E01013BF09404050F300",
INIT_06 => X"96F43FFF002004020044041084CB01AD000003761702401000FFDFE050000080",
INIT_07 => X"043C802A821D41412001A0040950AB60014114C3FE4187A009A663A680100B30",
INIT_08 => X"2C01004000047EFFF811A46968004060629A0002208A00000068113205A12034",
INIT_09 => X"0A812D8D5B742D3FF84056383FF7DE0880042107BFF9C45B85101C49A37F4000",
INIT_0A => X"0822189000480406310FFDFE00040009814C089202225412115414601DE3EBFE",
INIT_0B => X"C0281280080180B2948004400220011100841200D001000624000100C002804A",
INIT_0C => X"60694101816002D41A4068C101815004D8158809C86065941840B1014FFF56FF",
INIT_0D => X"0068C101816002D41A40694101815004D815810D42E04A08A80098C024500253",
INIT_0E => X"12682960828F05C96A001B029010134160C8125B0B271802242880A04482418A",
INIT_0F => X"100920C54E8EA256ECF078BA081C10080E05C0B06AA8B12CFD0D42E0441A3000",
INIT_10 => X"4F30A8801406D00290006280320100010362A8A20826A88660D86B202049F115",
INIT_11 => X"2011819E290048A2118EC8140C08064802C0081B0D64040936443306C5514410",
INIT_12 => X"C40A0300600C0A80509F418008804581BA0038005A706680012280506A801060",
INIT_13 => X"C000120080002341881F3FFFF80DCC158092C044600466208CC5091011C322A4",
INIT_14 => X"398C6021569249C4B3007127080806FF917FC30010107688862A28C54518DBFF",
INIT_15 => X"228D9228D9228D9228D99146C9146C84006309044081A001B188300E20806520",
INIT_16 => X"8004000000E07008010003EF80022A51904595123203040D9228D9228D9228D9",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010044800",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"0000000000004010040100401004010040100401004010040100401004010040",
INIT_1A => X"FFBFBFFF7CFE7F9E79E7FFEDDFEFFFBEFFE7DF83F7EFFFFDF7E0000000000000",
INIT_1B => X"FDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FBFDFEFF7FB",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800003FFFFFF",
INIT_1E => X"8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8001000040000000000",
INIT_1F => X"FFFFFFFFFFD74AA552E80010552EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A",
INIT_20 => X"2ABDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A800105D2EBFFFFFFFFFFFFFFFF",
INIT_21 => X"FFBD54BA552A800100000001FFFFFFFFFFFFFFFFFFFFFFFBD54BA5D2E8201000",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF7FBD74BA5D2E800BA5D00001FFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A552A800BA5D2E821FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E820BA5500001FF",
INIT_24 => X"FFFFFFFFFEFF7FFD74BA552E801FF002E975FFFFFFFFFFFFFFFFFFEFF7FBD74A",
INIT_25 => X"00008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA552A8200014003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E80",
INIT_27 => X"BDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2E800005D2ABFFFFFFFFFFFFFFFFFF",
INIT_28 => X"BD54BA552E82028002AB8FFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2A80000412A",
INIT_29 => X"FFFFFFFFFFFFFFEFF7FBD74BA5D2A800281C00001FFFFFFFFFFFFFFFFFFFFF7F",
INIT_2A => X"52A820AA490A071FFFFFFFFFFFFFFFFFFEFF7FBD74AA5D2E800AA5500021FFFF",
INIT_2B => X"FFFFFDFEFF7FFD54BA5D2E80082492E871FFFFFFFFFFFFFFFFDFEFF7FFD74AA5",
INIT_2C => X"0000038FFFFFFFFFFFFFFFBFDFEFFFFFD54BA5D2A801C7142E955FFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8000008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005D043FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"54BA552A80010002ABDFFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2E800005D2EBF",
INIT_30 => X"FFFFFFFFFFDFEFF7FBD74AA552E820BA002AA8BFFFFFFFFFFFFFFFFFFFFF7FBD",
INIT_31 => X"E800BA5D04021FFFFFFFFFFFFFFBFDFEFF7FFD74AA5D2A800BA5504021FFFFFF",
INIT_32 => X"FBFDFEFFFFBD54BA5D2A820AA082A955FFFFFFFFFFFFFFBFDFEFFFFFD54BA552",
INIT_33 => X"52E975FFFFFFFFFEFF7FBFDFFFFFFBD74AA5D2E80000082A955FFFFFFFFFFFF7",
INIT_34 => X"00000000000000000000002ABFFFFFFFFFEFF7FBFFFFFF7FBD74BA552A801455",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"8632CA211E4491D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"24B000808800040439245B221373581F97B0A8D1040F92000F42000047A00E58",
INIT_05 => X"011B2BBA308F023810004700083E220811E9BF2844021B1004045E4249500449",
INIT_06 => X"80A51003AA0200C020088E16A85235722940A817251101010100040D6D0702A2",
INIT_07 => X"5C9ECAB0D247B013B405EAD525FAE48FC2060B880081A26DCD4047EFF9EF0189",
INIT_08 => X"2D0141C0055280100751096B6A40D6F86723E510AA2004803D3275EB2024E814",
INIT_09 => X"04804818CD280100207246A8020000AC0283002004051507A5411C0DA0005048",
INIT_0A => X"2C6898B2950AA65635B00041C23020131A80CFDFF3FE509A907C556828201102",
INIT_0B => X"050F60E220A06880D2A14050A028501428054278142151262CA50343854E506A",
INIT_0C => X"612B3482C0C0078E1F412B1582C090078E1F840A2B0114020104022460002200",
INIT_0D => X"012B1582C0C0078E1F412B3482C090078E1F891C239F8908003099C1ACF06273",
INIT_0E => X"1BA859F213AFC14AA380430060181BA1B0FD16770236A4091621C08055C2C0DB",
INIT_0F => X"B08AA600CA88B143AB11880C280600101F09C030AB28B03C111C239F87082804",
INIT_10 => X"4B61BD8068B92400D0004E30368910E8822A984B0025B0DE6089462660095337",
INIT_11 => X"001AC2173B00E162563454C40804055412D4481128C4CC012A66F30455309600",
INIT_12 => X"50840180A00E1C81900C4190E160589C48082C006A9057CA4385809520F07830",
INIT_13 => X"004416B105036B4180C000800C8C00460848952220592745AC11A544B1BF0068",
INIT_14 => X"512C6A8C4F0008AA800470370000A0004D0000002126F30C902A29C54539C020",
INIT_15 => X"2A81C2A81C2A81C2A81C9540E1540E001400006100003202D040050220103D2A",
INIT_16 => X"22365034A8EA754008004C0214202C50013456520CA09281C2A81C2A81C2A81C",
INIT_17 => X"104411044110441104411044110441104411044110441104411044110445E220",
INIT_18 => X"0401004010040100401004010040100401004411044110441104411044110441",
INIT_19 => X"0003FFFFFFFF9004010040100401004010040100401004010040100401004010",
INIT_1A => X"FFBFAFBEFDFFBBBEFBEFBEFBDFD1FE3EFBD7ADF9B3EFDF7DF7D0512289000000",
INIT_1B => X"FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79EFFC",
INIT_1C => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000FE7F3F",
INIT_1E => X"8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2A8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8201008043FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74AA552E80010552EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E8000055",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD54AA5D2A82000552ABFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2A800005D2EBDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A800105D2EBFFFF",
INIT_24 => X"FFFFFFFFFFFFFFBD54BA5D2E82010002AA8BFFFFFFFFFFFFFFFFFFFFFFFFD54A",
INIT_25 => X"0100004000000000000000000000000000000000000000000000001FFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001008043FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74AA552E800105D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A820001400",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD54AA5D2E800005D2ABFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A80000412AB8FFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A82010552EBDFFFFF",
INIT_2B => X"FFFFFFFFFFFFBD54BA552E80038492EB8FFFFFFFFFFFFFFFFFFFFFFFFBD54AA5",
INIT_2C => X"00000001FFFFFFFFFFFFFFFFFFFFF7FBD54BA552E82028002AA8BFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201000040000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74AA552A820005D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001000043F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD54AA552E8001055003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"A820105D2ABDFFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2E800005D2EBDFFFFFFF",
INIT_32 => X"FFFFFFFF7FBD54BA552A80010002AA8BFFFFFFFFFFFFFFFFFFFFF7FBD54BA5D2",
INIT_33 => X"02AAABFFFFFFFFFFFFFFFFFFEFF7FBD74BA552E800AA082EA8BFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000000021FFFFFFFFFFFFFFFFDFEFF7FBD74AA552E820BA0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"5886C0201A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"0005EE040057700F40D08078500000D9218020407F0000BB8018A2FC380BEAC2",
INIT_05 => X"FFE0419028700023FCBC385F87C0BFFFE0124002FFE1E0C517FF09111212F300",
INIT_06 => X"16D03FFC96102081020000020489019C430480241202080810FFDFE000000000",
INIT_07 => X"0001160A003475C8100123400E20E1F40F439647FF4807E189A477EF81DF0AF1",
INIT_08 => X"801008000007FEFFFB110140695812CC4188D58A0AAA10803448D0844FB71000",
INIT_09 => X"4201258112D4487FF8001010FFF7DE4000000003BFF8C25818080020017F0F94",
INIT_0A => X"0C024000004A9400000FFDFF50010103134CAFDF03BA18000F39900037C3EBFD",
INIT_0B => X"C02812F00429DC92C40002000100008000105400C00400100000A01800080100",
INIT_0C => X"A1CAF13F214001521001CBF03F21100152100801C17E61841950B1C10FFF57FF",
INIT_0D => X"01CBF03F214001521001CAF13F2110015210088528E00E02C8200A430A424202",
INIT_0E => X"02C86040902AC60BACDF0E02D02001C1C044006D0C94FB94320880603C420B80",
INIT_0F => X"00010AF5052419D196441902801430182800A018D9CA8000648528E00D124802",
INIT_10 => X"4D101808458A5602E000892029110445C19960A00026880C006739000009B003",
INIT_11 => X"1009408021144CB042F880100C0601844068880CE72000013600600332C14000",
INIT_12 => X"F80E02120018390320F050144CB241D0B9023402085020825132C8CB5B404030",
INIT_13 => X"C200400020224000405F7FFFE0008E17C0D240406519400500840A9524EE38A1",
INIT_14 => X"AC810033149249C433200180082A06FF907FC308181204800600000000001BFF",
INIT_15 => X"010C1010C1010C1010C10086080860840063090442A18001B188300C48907120",
INIT_16 => X"0100000000000004002403EFC10302219A41C1443243050C1010C1010C1010C1",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200010",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000080200802008020080200802008020080200802008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000000000",
INIT_1E => X"8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8001000043FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2A8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA552A8200000043FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A552A8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8201008043FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74AA552E8000055003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2A8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E800000800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA552A8001008043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52A8200014003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8200008043FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74AA552E820101C003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E800105D043FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000043F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2A8001008043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"A8200008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001000043FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74AA552A820005D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552",
INIT_33 => X"5003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA552E8200055043FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA552E800105",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"0000745C200801000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"0001E6000053300F00D0007810042140C00000407F0000BB800000DC3801EA00",
INIT_05 => X"FFE0000008700003FC3C380F87C019FFE01240009BE1E00003BF00000000F300",
INIT_06 => X"06103FFC000000000000000004890088010080001202000000FFDFE000000000",
INIT_07 => X"0009B24B043980021000810284204A8001401643FE4007E5501AA00000DC8C30",
INIT_08 => X"0000000000007EFFFB11A56940581280031D61420000B080102040BC5B006120",
INIT_09 => X"020125811254083FF80000003FF7DE0000000003BFF8005800000000017F0000",
INIT_0A => X"0000000000000000000FFDFF4000000AA0354000019C40000128000011C3EBFC",
INIT_0B => X"C000104000000010440000000000000000001000C00000000000000240058000",
INIT_0C => X"4012500021B00880108012500021E00880104809C1666594584031010FFF56FF",
INIT_0D => X"0012500021B00880108012500021E0088010492064206100E81084200048C080",
INIT_0E => X"0410004C840041A0D8005410903804100144800803419043064900C002050184",
INIT_0F => X"020902F60002260D65B361BAA1041018140F02C0000809408D20642053027004",
INIT_10 => X"00020818B06D9802F00030C02060110002C9E8010C00010480B35A0300400041",
INIT_11 => X"20042108603100061516EE800C060228204300166B4060080008240593D00218",
INIT_12 => X"7C02000040206602C10B48110006143B62023C00142800B04400095DFF902030",
INIT_13 => X"C000000000000000001F17FFE000DC1180C7804400044029208301040214AE4C",
INIT_14 => X"008000010012414433000100080806FD107FC300000000000600000000001BFF",
INIT_15 => X"000C1000C1000C1000C100060800608400630104408180012188300C00814080",
INIT_16 => X"0000000000000000000003EF80020201904181003003000C1000C1000C1000C1",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"F30C2416857732AEBAEBFFA55EDCF9822659AE7BE742E6441990000000000000",
INIT_1B => X"3C1E0F07BEFBEFBEF9E79E79E79E79E7BEFBEFBEFBEFBEFBE7BE7BE7BE7BEC98",
INIT_1C => X"83C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F078",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8000001E0F07",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008040000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8001000043FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2A8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008040000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2A8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008040000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8000008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000043FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8000008043FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A800100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00004000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"4909E6093253306F82D0007C80000000080E01007F8020BBC00040DC3801EA00",
INIT_05 => X"FFE0000008704503FE3C380F87C019FFF01241009BE1E00203BF80800000F392",
INIT_06 => X"06103FFF9E2086C2086E006604C9019D03108B741202605040FFDFE070400880",
INIT_07 => X"4024057000000100000000000000000001401643FE4007C00000000000CC0830",
INIT_08 => X"0801404000007EFFFF40010000401408000045000000A0801000408000000000",
INIT_09 => X"4A7DF795965C6D3FFC0020003FF7DF01880C618FBFFDD75E00100040437F0000",
INIT_0A => X"0000000000009400000FFDFFC006020000000000019804000028000191C3EBFF",
INIT_0B => X"C02812E0182000F2C48304418220C11160845004D04820000000000000000000",
INIT_0C => X"0002400001000800000002400001000800000801C0786184185031810FFF56FF",
INIT_0D => X"0002400001000800000002400001000800000000202000000800000000080080",
INIT_0E => X"0000000404000000880000001000000001000000000090000008000000040000",
INIT_0F => X"000100C600800001040000040009100000000200200000400000202000020000",
INIT_10 => X"0002000000081001000000000040010000082000000001000001080000000040",
INIT_11 => X"0080000040010000001080001008000000010000210000000008000010400000",
INIT_12 => X"0000030280000000010000010000001020000000000000100400000108000040",
INIT_13 => X"E0120012C1400080291F17FFF0018C11808200400000400000C2000000042000",
INIT_14 => X"00800001001243443B000100880806FD107FC301800000000600000000001BFF",
INIT_15 => X"000C1000C1000C1000C10006080060840077330C4889CC292588300C00804000",
INIT_16 => X"82068C0200000008014023EF80020201904189003003000C1000C1000C1000C1",
INIT_17 => X"110441104411044110441104411044110441104411044110441104451044C820",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FFFFFFFFFFFFC110441104411044110441104411044110441104411044110441",
INIT_1A => X"200A625D144BC2B4D34D7F61432D518B45265EF8278C2015DA080800002FFFFF",
INIT_1B => X"88C4623124924924924924924924924904104104104104104124904124904281",
INIT_1C => X"58AC562B158AC562B158AC562B158AC562B158AC562B158AC56231188C462311",
INIT_1D => X"00000000000000000000000000000000000003FFFFFFFFFFFFFF800002C562B1",
INIT_1E => X"8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"0003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"94A7B2B1450000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"6FEBEF5FEC737AFBC6F85FDEB220109E1FEFFFE3FBA7FDFB9BD301DC3FF5F0D2",
INIT_05 => X"FEEDBFDC387F987FEF7C3FAF87FF59F7F5FB7FF59BE1FF980BBBB7FE6D21F3DB",
INIT_06 => X"57902FFDEE9D7DC9D7DF2B263893479DDFAFDFE15213FEFEBFFFFBE1F1D3A333",
INIT_07 => X"10992310605CE10301DE0C1831CB7DF60A244B9BFEE00589DDBCEFEDC1DFA089",
INIT_08 => X"001D8EA111DA7FEFF90F21C8C84D9C0D858FC7020828C18FD18346BBF0000180",
INIT_09 => X"F37DF7B9DF7DCB3FDE89ECC07DF7DF5F985C6BCFFBFA28F99E7EB07F47FFEFAA",
INIT_0A => X"7DCFE1D4077B4D0026FFFFBE7D67D7F3BB79CFFB83BF14EC1E7D5980580BFAFF",
INIT_0B => X"C7D7D51D6F5FDCB935D7AFEBD7F5EBFBF7FEBD66DBFCA3F87501AE7B08060730",
INIT_0C => X"01F45EC0010007E01001F45EC0010007E010084BCD7FF1B61B5C33813FFFFCFF",
INIT_0D => X"01F45EC0010007E01001F45EC0010007E01001BD8020500008001F0100405202",
INIT_0E => X"1EC00040B02007EC09A0E00010001DC0004600400F781429C0080000770001A0",
INIT_0F => X"404B3BFD0402346235408402C08010003C064000E408010081BD802060020000",
INIT_10 => X"0E401A08FE0012040000FC002001360403E434588007200D00F88C84C081C203",
INIT_11 => X"001F01002156040675809145400007B00040091F1190982038406807C868B100",
INIT_12 => X"008320C0403C34000088601604067D00212000007C400082D81009FC08281D00",
INIT_13 => X"F7BFFED3FBFF6A84383F177FF005FFBFF5FA1040076065F730FC08043A903A80",
INIT_14 => X"F589807B7096CD4CF73AC1FC98884FFF19FFC71FEFED7B251E35768E8ED6BFDF",
INIT_15 => X"8C0D78C0D78C0D78C0D7A606BC606B8C56F7730ECCDBDF152199F51EDDCDEBCF",
INIT_16 => X"DFE7DD87FEFF7FF796FFFFFDFFD7E681B867D3683A03A40F78C0D78C0D78C0D7",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFEFDFD",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"FFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEB",
INIT_1A => X"57AA9ABAD8ACBF0E38E3A89F9E923C2CD990A7D0D2A377F86EDB5C88646FFFFF",
INIT_1B => X"4C261309861861861861861861861861861861861861861861A69A6986186EBC",
INIT_1C => X"84C26130984C26130984C26130984C26130984C26130984C26130984C2613098",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000261309",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"1085B0B041000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"6FAB975B6470BAF386C87A9CB00000001FEF9F23E3A7BDE79B5101D23FB5C0C2",
INIT_05 => X"F8EDBFD4347F18778E723F2E47FE59C7F5FB7F759B91FB880BA3B6FE2921CBDB",
INIT_06 => X"47000FFC128D5CE8D5CC210638A046889CAB57E8421786B6ACFFE3E181932377",
INIT_07 => X"000000042000000288020C18300320620A80231BFE200181092CE7ED80DFC001",
INIT_08 => X"000C562551D87E8FF90041101042110180004102800008801183468180000141",
INIT_09 => X"137FF7A0FF75813F1C85244071EFBF17D85C738BE3FA08F9DE36B05B07FEEF22",
INIT_0A => X"768EA0C406630D00226FFE3E2D62D6E21259CFDB039E806C02451880400BE0FC",
INIT_0B => X"CC57550D63564D1D2556ADAB56D5AB6AD7EAB962CBD8A3A83101F47E08040510",
INIT_0C => X"01E44A40010007600005E44A4001000760000843C561E5C55C42B9011FFF48FF",
INIT_0D => X"05E44A40010007600005E44A40010007600004BD8020100008001F0100001302",
INIT_0E => X"1EC00000382006EC0820A00010001DC0000208400D781020C008000077000020",
INIT_0F => X"40431BC50402146235400400408010003C064000C400018080BD802020020000",
INIT_10 => X"0E400204FE0010040000FC0000003E0403A424108007200102E888808081C200",
INIT_11 => X"001F0100005E040475808101400007B00000015D111010203840081748482100",
INIT_12 => X"00012040403C34000080201E04047D00202000007C400000F81001FC08080500",
INIT_13 => X"E5ADA4C25ADE72041A3F147FF0018DBBB5FA10400360649310FC08003A903A80",
INIT_14 => X"054880693016DD4C755AC16C1A884FFE18FFD757E7ED7A211E81C09818109E1F",
INIT_15 => X"440C3440C3440C3440C3C2061A2061AD46FF730E5CCBCD55219AB55F0DEFABC7",
INIT_16 => X"5EC71385FC2512E3565BBBF1BAD6F281BC63F1683803C00E3440C3440C3440C3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BDE75ED",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"FFFFFFFFFFFFAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB",
INIT_1A => X"200E5E48710A4200000028150200903950C086D0E28028104A471688747FFFFF",
INIT_1B => X"0080402000000000000000000000000000000000000000020800000000000780",
INIT_1C => X"5028140A05028140A05028140A05028140A05028140A05028140201008040201",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8000028140A0",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"8C2100804900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"02000100440408002408008002221000204116A280000F000001400000100010",
INIT_05 => X"0004D44400004D4400000000000000000000005C0000000A0000002C20600000",
INIT_06 => X"4100000120040A0040A00B0090006202940100004000A2020400200888800911",
INIT_07 => X"5002489020420110800244891211440804000810002000081040000000200000",
INIT_08 => X"080542C004CA00000050080202008401842004108AAAA00008912240A1248804",
INIT_09 => X"0000000C0000E400002040500000009202C1002040004400022200020400B062",
INIT_0A => X"58C460540329810002D002000400407020800000004000640800088008280001",
INIT_0B => X"0140000401028008330000800040002002480102010082981500062108020430",
INIT_0C => X"00040A40000000A00000040A40000000A0000040060084104110828030000800",
INIT_0D => X"00040A40000000A00000040A40000000A0000000800010000000000000005000",
INIT_0E => X"00000000A00000040020A000000000000006000000080020C000000000000120",
INIT_0F => X"4040152000000020000004004080000000000000240000000000800020000000",
INIT_10 => X"0000120002000004000000000001220000040410800000090000808080800002",
INIT_11 => X"0000000001420000200001014000000000000900101010200000480008082100",
INIT_12 => X"0001204000000000000820020000200000200000000000028800002000080500",
INIT_13 => X"00933050080C0001900020000000408010000000022000D61028000008000000",
INIT_14 => X"400082D022040000400800081022C0000080000206CB0821082B694D4D294000",
INIT_15 => X"050160501605016050160280B0280B0012000843066021001400040024440245",
INIT_16 => X"0861CD33548542A10209D4100E4040A00002002C004001036050160501605016",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008021081084",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"0000000000000020080200802008020080200802008020080200802008020080",
INIT_1A => X"06A0A0F108816B1861863BED822140048D2E5818732C5589A40A0C22E1000000",
INIT_1B => X"80C0603020820820820820820820820820820820820820820820820820820035",
INIT_1C => X"582C160B0582C160B0582C160B0582C160B0582C160B0582C16030180C060301",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800002C160B0",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0803B2814D0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"26E1E905CC574828C4F85FC600000016004F77E2F887CDB80BC340DC07D1F000",
INIT_05 => X"FE1DFE4C080F884FE33C078F803F19F011E93ED49BE01F1A03B8972E6D20F049",
INIT_06 => X"57902000DE142D4142D5030010134395D70589415002DA4A17FFF800F0C38111",
INIT_07 => X"00092300601CE00101DE040811D919F402244293FEE00400CCB46BA4C164A088",
INIT_08 => X"08148A4000887FE0000F20C8C80D080D818FC2000000418FD08142BAD0000884",
INIT_09 => X"E204D2154D28AA3FC60888D03C10415A80402847F8002458926A002E457FA0AA",
INIT_0A => X"5587A1540231410006DFFF80540541619968C76980E914E4163D4980100BFA02",
INIT_0B => X"07C7C0140D0B50A8218102C0816040B1225C1506512C83E85500AC3A08040630",
INIT_0C => X"00141EC0000000A01000141EC0000000A01008480D3EB4A24A0C910037FFFC00",
INIT_0D => X"00141EC0000000A01000141EC0000000A0100100800050000000000000405200",
INIT_0E => X"00000040B000010401A0E000000000000046000002080429C0000000000001A0",
INIT_0F => X"40483B590000202000008402C080000000000000240801000100800060000000",
INIT_10 => X"00001A08020002040000000020013600004414588000000D00108484C0800003",
INIT_11 => X"000000002156000220001145400000000040090210909820000068008828B100",
INIT_12 => X"008320C00000000000086016000220000120000000000082D800082000281D00",
INIT_13 => X"32936E43A92F2880B01F37001004B29450580000066021F6303C000408000000",
INIT_14 => X"B481806A62840800C22800B8900042FF0180000ABFEF89250815568A8AD6ABC0",
INIT_15 => X"8D0068D0068D0068D006A68034680300021410028450530014014002D445624D",
INIT_16 => X"89418D13FE7F3FFD8BADB7FC4F4164A00806522C0A40A50268D0068D0068D006",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C4B12C9894",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"FFFFFFFFFFFFC0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0",
INIT_1A => X"FFBF3F5E7CFC7DFFFFFFD7FADDCFFFBEFFCF1F879DFFFFFDFFEA0C00602FFFFF",
INIT_1B => X"DFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBAEBAEBAEBAEBAFFFD",
INIT_1C => X"FDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800003EFF7FB",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"F7AEBEBFFDFFBFBEFBEFFFFFDFF3FC3EFFF7FDFBF76FF7FDFFD0000000000000",
INIT_1B => X"FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79EEBD",
INIT_1C => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000FE7F3F",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"1084B030000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"6DA986092050306382C05A1C900000001FAE89016387B2A38B5000D03FA1C0C2",
INIT_05 => X"F8F92B90307F41338E303F0E07FE19C7F1FB7F289B81FB8003A396D20940C3DB",
INIT_06 => X"06000FFC020004C0004C000628800488080003600213001000FFC3E101030222",
INIT_07 => X"000000000000000220000810200220620E00030BFE000181092CE7ED80DF8001",
INIT_08 => X"0000000001107E8FF90001000040100000004102200000801102448100000100",
INIT_09 => X"027DF780DF74013F1C00240071E79F05888C618BA3F800599C101049037E4F40",
INIT_0A => X"240A808004420400202FFC3E002202021259CFDB039E0008024510000023E0FC",
INIT_0B => X"C407500020004C10060204010200810040801060C04821202001A05A00040100",
INIT_0C => X"01E04000010007400001E0400001000740000803C0616184184031010FFF40FF",
INIT_0D => X"01E04000010007400001E04000010007400000BD0020000008001F0100000202",
INIT_0E => X"1EC00000102006E80800000010001DC0000000400D7010000008000077000000",
INIT_0F => X"000308C50402144235400000000010003C064000C000010080BD002000020000",
INIT_10 => X"0E400000FC0010000000FC000000140403A020000007200000E808000001C200",
INIT_11 => X"001F01000014040455808000000007B00000001D010000003840000740400000",
INIT_12 => X"00000000403C34000080001404045D00200000007C400000501001DC08000000",
INIT_13 => X"E004048240426200081F147FF0018C1380DA10400140640100D4080032903A80",
INIT_14 => X"050800A91012494C31004124080886FE187FC301B124F2001600000000001A1F",
INIT_15 => X"000C1000C1000C1000C18006080060840477330C4889CC012188310E08812982",
INIT_16 => X"02061004A820104809402BE1900222019861D1403803800C1000C1000C1000C1",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100446020",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"FFFFFFFFFFFF8100401004010040100401004010040100401004010040100401",
INIT_1A => X"00000000000000000000000000000000000000000000000000001000802FFFFF",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000000000",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"88280C4C7B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"00160090920C04800904848262220277E05152B280780D407428E723C01E1400",
INIT_05 => X"0006D46207801E400183C0707800E6000E008057641E00473C40680D32330C00",
INIT_06 => X"C165000225E2C11E2C12A0D0144AC27206582C166504816162002000B0FC21D5",
INIT_07 => X"5E6D233B964E7CD99DFB870E1DDDD889C5FBDC440129A0604442180238203F70",
INIT_08 => X"AD23C17544C581000657A0E8E83D86F0E4A7B2D88AAAFD7FE0E1833AC5920CFC",
INIT_09 => X"6D82082E2081B6C0027ADA398000008A504318404005B70663212C04A080B036",
INIT_0A => X"414568729139FA5610C00001A2502440888420247041E87681008CE9AFC80001",
INIT_0B => X"22B826E250B12346F1244812240912048941621804A150CA1CA45C254D4AF4AA",
INIT_0C => X"F80FA97FE0F0009E0FC40FA97FE0F0009E0FC048211E9C11C31F82E4A0008900",
INIT_0D => X"040FAB3FE0F0009E0FC40FAB3FE0F0009E0FCC42EFDFBF0AE03080E2AEB2E0F1",
INIT_0E => X"013879BA878FE807F65FBF12E0380231F0BD9E3FC08FEBD6F661C0E008C3CB5F",
INIT_0F => X"B248831ACBFC8BBDCAB779BC699F20180309A0F83BE2B87C7C42EFDFBF187806",
INIT_10 => X"4131B59003FFEC07F00003F01FB90BE9F01FC8B38C2098DAE007F323A0C83136",
INIT_11 => X"3080E29F1B2BE9F8A27E6E915C0E004C72BEC800FE7464290626D7003F994718",
INIT_12 => X"FC0C2352A0024B83F07F198BE9F8A0FFDA2A3C0202B8776A2FA7F023F7D06570",
INIT_13 => X"1448126105810941C5C068000CD4004C0905E52630BB1AE49C2BA7F98D6F846D",
INIT_14 => X"6074EA560F0416A24844B01302A26100C4801844069B0C88881A28C141118000",
INIT_15 => X"A781E2781EA781E2781C33C0613C0E21020800239450116ED443C041B47E9665",
INIT_16 => X"241140A056954AB0C280D0002020187007122C3E04E03383E2781EA781E2781E",
INIT_17 => X"20481204812048120481204812048120481204812048120481204812058112C1",
INIT_18 => X"0481204812048120481204812048120481204812048120481204812048120481",
INIT_19 => X"0000000000001204812048120481204812048120481204812048120481204812",
INIT_1A => X"C4109CAF9C4C83B8E38E2AE9C136AD8E9B562CF042E6281CF13043A85D400000",
INIT_1B => X"F0F87C3E08208208208208208208208208208208208208208208208208208220",
INIT_1C => X"1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1",
INIT_1D => X"000000000000000000000000000000000000C3007FFFFFFFFFFFA00000F87C3E",
INIT_1E => X"4214555517DEAA5D7BFFEAAF7803FEBAF7FFD74BAAAAABDEBAF7AE8000000000",
INIT_1F => X"1555FF55517FE000055421FF00557DF45A2D5401EFF7D142145A2AE800BA0851",
INIT_20 => X"5555555A2AABFFFF5D516AA00A28028A00AAAEBFE00A2FBD75FFFF8400155085",
INIT_21 => X"5517FF45A2AEBDEBAAAAAA8BFFF7D140010FF84174BA552EBDFFF0004020005D",
INIT_22 => X"5504000BA5D2E97545A28028B4508554014508043FEBA082ABFE10AAAEA8ABA5",
INIT_23 => X"FA2AABFE00FFFFD74AA085540000002E801FF557FD75FF0051401FF5D0015410",
INIT_24 => X"EFF7FFC20BAF7D1575450800020BA08517FF45F7FBFFF45A2FFFDE00002E801F",
INIT_25 => X"A38BF8FC000000000000000000000000000000000000000000002ABEFAA80001",
INIT_26 => X"7155BC2A87092AAFA9257F1C5BC00AA5D7FF8EAA57803AEBAF7F5D74AAA2A03A",
INIT_27 => X"BFBC7EB8005B55A85B555EF095F50578085BE8FC7A3F00516DA2D5451D7EBDB4",
INIT_28 => X"0975FFAAA1521FF492BF8F40B6AAB84AF555168A00EA8000150A801C01C7142E",
INIT_29 => X"2EBAE28168ABAA2D43D568BC5400168E90E2F412BEAE3D542A004380124921D2",
INIT_2A => X"2FA3AA28EA8168A954100071D2E90A855C7A00A38F6DE05B40480557A95A3A1C",
INIT_2B => X"16D1EAE925EA0BFEBF4AA09217F490568417085147B50A80095178157FEFA074",
INIT_2C => X"000002D57AAA8402A8743DBD202DA95568A95E800A8F57F6DA971F8F7FFFA42D",
INIT_2D => X"AAFFD1564BA2282BFA02A2C28000000000000000000000000000000000000000",
INIT_2E => X"5EFA87F57555AAFBD7555FFAE95408A8FDC31AD017D34ABA5D7BEAAAAD786BCE",
INIT_2F => X"C2087383F79A5046A37B55F38415555797D63BFF007F8B2B2D97D483AFA7BD9F",
INIT_30 => X"42000D382964A92B401E71D7581C33172EC0A0300A6AEA8FAF0451CA001D4845",
INIT_31 => X"C8365A2FD5E04AA5780A8AAAD7AC3CA02003BEBBA7D7463CC508D07577BAFBD5",
INIT_32 => X"0621F562B1122DA70C3808458881056A5502AA150502828811FCD4EABDB1DFDF",
INIT_33 => X"96D55BBAAC55EAFAF86D35E4A92B4460D15060374FF72AAADF24559515705079",
INIT_34 => X"007FC0000007FC0000007FC07AAF12E00505D3FDF6A03D4BFB79AFA4C5CB5F58",
INIT_35 => X"0007FC0000007FC0000007FC0000007FC0000007FC0000007FC0000007FC0000",
INIT_36 => X"00000000000000000000000000000000000000007FC0000007FC0000007FC000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000040000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"CA1800080848B0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000010822C00803804000001999EF9C00040B0002000001000640200001018",
INIT_05 => X"0000400244000000014200004000000004000000001000032000200002100800",
INIT_06 => X"208500000080412804100CB08000302220080408010000202000000404100844",
INIT_07 => X"5AF6FEF002230018010860C1833C460044204C000008A0041000080008202800",
INIT_08 => X"8D22C0F55000010000524481890BC000263000188AAAA10F8C1830562B25FC4C",
INIT_09 => X"B102002E20013600022D8819000000A000110A4000002C204000240420001000",
INIT_0A => X"02605C1C1108481200C000002040040820000020104100028800002801041001",
INIT_0B => X"081001004010810510040802040102008100200800A1100707040101E20BE0B0",
INIT_0C => X"58000003C0F000A000C4000003C0F000A000C0000012187087010AE4B0000000",
INIT_0D => X"04000003C0F000A000C4000003C0F000A000CC4200002F08E03080000010F180",
INIT_0E => X"0000000AAC00680000001F10E038000000078808C00000023461C0E000000127",
INIT_0F => X"5200040A00D000000202090C281F201803000000240218C0044200001E187806",
INIT_10 => X"400012900001EC03F000000000392100B00048230C200009A000130320480002",
INIT_11 => X"308000000961002880204A901C0E00000002C9000260640900004D0000904618",
INIT_12 => X"5C0C0312A002000000083881002880025A0A3C020000002A8400B00007806070",
INIT_13 => X"04080830008010468220A00008D0000801046004308A18500002012800090428",
INIT_14 => X"0840280206089000004090110200000000001454000200828008081110084000",
INIT_15 => X"4191AC191AC191A4191A00C8560C8D2910000060901010401E13405111220000",
INIT_16 => X"0410028000100800140000002004103224002006406401918C191AC191A4191A",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200800041",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"0000000000000200802008020080200802008020080200802008020080200802",
INIT_1A => X"2431A589945201924924B060D757DF8A94102E038728287452B4008A04000000",
INIT_1B => X"75BADD6EAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8A28A28A28A28AB20",
INIT_1C => X"974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D6EB75BADD6EB",
INIT_1D => X"00000000000000000000000000000000000303FFFFFFFFFFFFFFC00000BA5D2E",
INIT_1E => X"FDFFFA2FFD74000855555FFFFFFC01FF087BE8BFF5D2AAAB5555554000000000",
INIT_1F => X"EBFF455D04175FF5D7FEAAAA002ABDEAA5D2EBFFEFA2D17DEBAF7D1574BAAAFB",
INIT_20 => X"8415400005540155F7D16AB45002EA8ABA005540145557BFDEAA5500154AAAAA",
INIT_21 => X"5003DE00A2FFFFFEFAAD57DE00082AAAA00082A820BAAAD540145F7D5574BAAA",
INIT_22 => X"F7D5554AA5D2ABDEBA082A821455D2EA8B455D2A975EFF7AEBFF550055555FF5",
INIT_23 => X"FFF84155FFFFFFFFF55AAAABFFFF5D556AB45A2D16AABAAAAEBFE10AAFBD7545",
INIT_24 => X"10FF84174BA552EBDEBA0004020AA5D04155FFAAFFEABEFA2FBEAB455D7BD55F",
INIT_25 => X"F47015A800000000000000000000000000000000000000000000175FFF7D1400",
INIT_26 => X"FEAAF7D5524AAA2F0BAF7FABDFC7E10005F525D74BFBC51FF1471E8BEF55242F",
INIT_27 => X"50492490E17EAAA2AAB8F4515043DFC75575C7000B6AEBAEAA5D2EBDFFFBED17",
INIT_28 => X"B6FB6DF7DFD5038ABA140A2D00554517DEBDB6FB55142A8708202FBD257F1C75",
INIT_29 => X"AABFF55BC5B555C74B8A38E38085BE8B47A3A00503D1420AD000B420820AAE2D",
INIT_2A => X"AABD21EF1C2FEA5FDEBDB505FA4920AFE10082E925555F8FFDE38087FC51C7F7",
INIT_2B => X"1EFBFDBFF5FF1C00BF5D25475C7B7FEAFF45BEAABA4AF555168B68FEDF6AB52A",
INIT_2C => X"00000151EAE3D542A004380124921D20BFFFA0AA17AEB8BFF155552B6F5E8BFF",
INIT_2D => X"FF55516ABEFDD003EFE5093DC000000000000000000000000000000000000000",
INIT_2E => X"2BA5D2ABDFFFF7D57DEAAFFD5420B2A2D37DB07A3D795000087BC01458AFBC11",
INIT_2F => X"D608897FD610D01151C610592A974BAFBAC28B55550434D555C53E0CE2AAA874",
INIT_30 => X"3FE102400144ABAAFFF7DE772FDD56588042F72EF0851575FFAAFBDD5542B2ED",
INIT_31 => X"F6A81A239501755F504BDF557D79431FD006EABA100F3D68FFFAABAC20EF0400",
INIT_32 => X"55EAF57FF957CAAA7FABF7DFD0C6A7DFFFA07FC04EA0006BFE007E2E8315DD02",
INIT_33 => X"FADF6900FFFF68BEFDFFB4B1FE5551141E78A02803158517BD745AEAEA8FAF0C",
INIT_34 => X"0000000000000000000000165BAFBD542000D382964A92B403EE18D5408A6F2A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000040000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0812",
INIT_01 => X"A145A00810790848048044A54E404340404000720885800802000906E4910200",
INIT_02 => X"5C010802020408040C455850AA055254090541A111200A104A0000000908B510",
INIT_03 => X"182002200C00004485264A001214912802150020218808002440854288890550",
INIT_04 => X"210302008014100120806B08702010102722C9E0412200651102418214049492",
INIT_05 => X"48416A98042912208552102442884882A58A08011290A1120A81230240018DCA",
INIT_06 => X"12800554528021C8023A28000031240048000100001170000155414109102066",
INIT_07 => X"000022104040810089080810211A04480420420154800088096A0EA8C0222080",
INIT_08 => X"080198C105424705510A08828A0B19080428040080A0A10F8102049300000804",
INIT_09 => X"3165541CD54822160A89E89020AA8AC4CA1D39CE215264B04040002400B80688",
INIT_0A => X"280201840548C80001C568146000001012D40D7182411080153801004800B057",
INIT_0B => X"4812050000080114100206000100818100900640C04C20104101021C00000310",
INIT_0C => X"00A00000010000A01001400000010000A0100801407234E34C1A980001552055",
INIT_0D => X"01400000010000A01000A00000010000A0100038000000000800000000405000",
INIT_0E => X"00000040A00002600000000010000000004608000850000000080000000001A0",
INIT_0F => X"400020C4000200420040000000001000000000002408000000A1000000020000",
INIT_10 => X"00001A04940000000000000020012800018000000000000D0288000000000003",
INIT_11 => X"0000000021480000508000000000000000400951000000000000681300000000",
INIT_12 => X"00000000000000000008600800004C000000000000000082A000015000000000",
INIT_13 => X"80004012C06000018004342AA000700000000000044000500000000022101800",
INIT_14 => X"958100134200904487400010022005E0110D524029263100009200151409130A",
INIT_15 => X"C9013C9011C90134901144801A4808AD4451394CD0391A541593C04B59084008",
INIT_16 => X"010400A0A890684444240120C0071420344423040240450114901149013C9011",
INIT_17 => X"080601806018060180200802008020080601806018060180200802048026C000",
INIT_18 => X"8000080001804018040180400800008000080601806018060180200802008020",
INIT_19 => X"1F83F03F03F00180401804018040080000800008000180401804018040080000",
INIT_1A => X"E90C042CB002102CB2CB2EE00271AE180616A85246C77250C7D00022012F81F8",
INIT_1B => X"28944A2504104104104104104104104104104104104104104104104104104608",
INIT_1C => X"128944A25128944A25128944A25128944A25128944A25128944A25128944A251",
INIT_1D => X"000000000000000000000000000000000003C3007FFFFFFFFFFFCE3F00944A25",
INIT_1E => X"EAA1055042AA105555421EFFFD568AAA002EBFEBA550002000AA800000000000",
INIT_1F => X"AA8BEFAAAE975FFA2D5555450851574000851554BAFFAE801FF087BE8BFF5D7B",
INIT_20 => X"2EA8AAA5D2EBFFFFA2D1554BAF7D17FEBAAAFFFDFFFA2D57DE10557BE8ABAF7A",
INIT_21 => X"D04175FFFFD5574AAAAAA974BA082EA8BEFAAD555555F7D568ABAF7D5574BA55",
INIT_22 => X"085557410F7AA97410087BD55FF087FEAA10A2FFEAAAA552AAAAAAAAAABFF455",
INIT_23 => X"05D7FE8B45F7FBFDE00085540155F7D56AA00007FEAA000055401555D7BFFE10",
INIT_24 => X"00082A820BAAAD540145F7D557410AA8428A10550017400550402155A2803FE0",
INIT_25 => X"000E28A80000000000000000000000000000000000000000000017400082AAAA",
INIT_26 => X"01FF1471E8BEF5574AFA00010ABFA38555F401D74BD16FAAA002ABFEAA550E82",
INIT_27 => X"FF400417FEF082F7AAA8BEFE2AA955EFA2DB5757FEAFBD2410005F57482E3AA8",
INIT_28 => X"F6DA82F7DF520385D2FE80AA5D2EBDFD7BED1574AAF7D5524AAA2F1FAF7FABFB",
INIT_29 => X"24ADAAAB6AAB8F455784155C75575C7000B6AE95492082EADBFFBEDB55555E3D",
INIT_2A => X"051C05571474024A81C5557578EBA087400007FC21C7005B6FB47F7A438E925D",
INIT_2B => X"E10A001FFB40038F68F7F578F7FFEF568E2808554717DEBDB6FA3D0075EDA800",
INIT_2C => X"000001043D1420AD000B420820AAE2DB4716DF7DFFDE381D716FA15550015428",
INIT_2D => X"AA002ABDEAA552A80010AAA88000000000000000000000000000000000000000",
INIT_2E => X"800087BD5410AAAA801FF55556ABEF5D517EEE00828FDEBA5D7BC015582D57DE",
INIT_2F => X"A2B2A3D169B07A3D7BFE10597BFDE00AEAC28BFFAAAE955EFAAFBC15F5A3D7D6",
INIT_30 => X"BDFEFFFFBC1154AAFFFFE107FF9D72A20842080BA5D2ABDF55F7D575EAAFFD50",
INIT_31 => X"97CF4780286A2105D2A3FEBAFFAC28B555504145555A53C00B2A2AA02000082A",
INIT_32 => X"FFFDA02003FFDEAA8557D65550915544AA5D51574EAA28015400547FC315D007",
INIT_33 => X"16F9E2555500174AA282E20BFFFF842AAAAADD5699ADABD5A8AAA0051575FFA2",
INIT_34 => X"0000000000000000000000030EF04003FE102400144ABAAFFD75E7F2BDDD2B80",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000080000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380202",
INIT_01 => X"200C9A424080216D3C2462C99E104B49404040028804A0080A000416A8D90A0C",
INIT_02 => X"4809A902031800444461089C66E331352180D468B8240E600C0081110B80ACD0",
INIT_03 => X"DA16C2210C0001D231A30A0648C68428320066010A80881068A80C401CC46330",
INIT_04 => X"2088601DA82700EC92307064A3756910088469A01C250210990240420E005A48",
INIT_05 => X"2D2060182414411A314A0A02C18C01B9854368080A506912018C2502484038D1",
INIT_06 => X"16801CCCAA8061E8061C0D008020140520080769000420202133CCC50C110804",
INIT_07 => X"5800B65040630008810C20508138071604A461833280038C89904E6400232008",
INIT_08 => X"0800906010521D1CC80204918949540C061000088000A90F840A50963A017845",
INIT_09 => X"A037A02C68552A35620C88900A69876100810A6A84C82C400040300D40D20A48",
INIT_0A => X"062A10B40042C80000CCE4CC2045051913208CE80243048008204100402079CC",
INIT_0B => X"C81301004C18912102060C0207010201C190200400A401042D00F15884030170",
INIT_0C => X"0190148000000800100450148000000800100401CB33494594532980733322CC",
INIT_0D => X"05101480000008001004F014800000080010051C000040000000000000480000",
INIT_0E => X"00000044000001680180400000000000014000000B1004090000000000040080",
INIT_0F => X"00812E44000024400140800280000000000002000008000001B0000040000000",
INIT_10 => X"0002080CCC0002000000000020401000034010480000010402D8040440000041",
INIT_11 => X"00000000601000064180104400000000004100570080880000082015C0209000",
INIT_12 => X"00820080000000000100401000061C0001000000000000904000094C00201800",
INIT_13 => X"4408400000A26285A03224E670094008010000004444010E2050000420801880",
INIT_14 => X"4DC10283429294408740C0B48202854C011CD75C0102A30400A8891451284B26",
INIT_15 => X"4901A4901849018C901A648056480C2D4449116DC0115C41159B655F112AC008",
INIT_16 => X"0510000000DA690C1D20030BA0011421B404220402404501A49018490184901A",
INIT_17 => X"280803808038080380803808038080380C0280C0280C0280C0280C0680C28051",
INIT_18 => X"00C0280E030080380A030080380A030080380C0280C0280C0280C0280C0280C0",
INIT_19 => X"B556AA9556AA830080380A030080380A030080380A0200C0280E0200C0280E02",
INIT_1A => X"742C000A981E80249249206018F18E0C85142822266800586291000A844D54AA",
INIT_1B => X"A9D4EA7524924924924924924924924924924924924924904104104104104A20",
INIT_1C => X"1A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A753A9D4EA753",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF849010D46A35",
INIT_1E => X"42000AA802AA10F7D57FEAA557BE8B45A2D5555EFAA800015508000000000000",
INIT_1F => X"BC0155A280021EFA2FFE8B4555042AA105555421EFFFD568AAA002EBFEBA5551",
INIT_20 => X"D5574000851554AAFFAE801FF087BC01FF5D7FEAA10550402000AAD56AAAA557",
INIT_21 => X"AAE975FF005540145A2D157410AAD17DFFF5D0400010AA842AAAAFFD542000FF",
INIT_22 => X"F7AE975FF080428B455D7FFDEAA5D55574BA00517DE105551420BAF7AAA8BEFA",
INIT_23 => X"F007FFFEAAAAD5554AA552EBFFFFA2D5554BAF7803DEBAAAFFFDFEFAAD57DEAA",
INIT_24 => X"EFAAD555555F7D568ABAF7D5574BA552E800BAAAAE800AA087BD5555552A821E",
INIT_25 => X"155080E800000000000000000000000000000000000000000000020BA082EA8B",
INIT_26 => X"FAAA002ABFEAA555E02000E28AA8A38EBD578E82E975EAB6DBEDF575FFAA8E02",
INIT_27 => X"87A38AAD56DA824975C217DAA84021FFAAF5EAB55EBAEADA38555F451D7EBD16",
INIT_28 => X"E2DABAFFDB47412ABFE90410005F57482E3AA801FF1471E8BEF5575EFA00012A",
INIT_29 => X"5F47082E3AAA8BEFA02A955EFA2DB5757FEAFBD2400BED57FFD7410E05038BE8",
INIT_2A => X"2F1FAF7FABFBEAE2AEBA4974871C043AB6D4975FFEBA5D71D742A407FFFE0055",
INIT_2B => X"1C75D25C74920821D708757AE2AA3FFC04AA552EBFFD7BED157482F7803AEAAA",
INIT_2C => X"0000007092082EADBFFBEDB55555E3DF6DA82F7DF7AE38497FC00BAB6A485082",
INIT_2D => X"FFFFFFD75FFAAAE8014500288000000000000000000000000000000000000000",
INIT_2E => X"EBA5D7BD5545A2D57DEAA002EBDEAA557BC0010AAA8A8ABAAAD568A1020516AB",
INIT_2F => X"29EF5C517EEE00828D74AAFBD57DE000057C21FFAA80001FFAAD57EB55A2A8AB",
INIT_30 => X"7DF55082E974AAFFAABDEBA77FDD66A0ABBDC2000087BD5410AAAA801FF55556",
INIT_31 => X"7C14100957FF6105D7BD5400AAAC28BFFAAAE955EFA8FBC15E5A3D5D7400FFD5",
INIT_32 => X"D1554A8FFC42AA10A7D169F57ABD7FEEBAAA841550555002ABFF54517EEB25D5",
INIT_33 => X"96F014AAFF84154105555C215500000014558557FA42A3D7020BA5D2ABDF55F7",
INIT_34 => X"000000000000000000000015400082ABDFEFFFFBC1154AAFFFFE10FFF9DF2020",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000040000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204002",
INIT_01 => X"010398000008004C1C20650E1E104348403008418984014902030006A0910200",
INIT_02 => X"480108A200000000444048E41E80F00A4104311868200200080000000988A390",
INIT_03 => X"0CA08220080000D004060A0240101028270012603000000030808C0208C000F0",
INIT_04 => X"4403A609A055306BC2C0735810CEE5100A0A40E06B8360E3808241D03845D002",
INIT_05 => X"ECE0498800791403AD3038AE079059A790E245819A41E4120BAB87800001D312",
INIT_06 => X"06000C3D220003E0001A210088B1008C4004034912120000010FC3C00000A064",
INIT_07 => X"5000220440000000090800002118400204206100F040018019004B8001232088",
INIT_08 => X"0810884441123323C0424180880B0108002000000880890F9000041200000845",
INIT_09 => X"230B6715A4786E0F5A8C889031EF9F45D884794FA03A24781840100D000E1140",
INIT_0A => X"0C4202200142400004DC3C82600401003200872003FB1400082840001022003C",
INIT_0B => X"C800940008088034040000010000808140901000C00001008800A01814000840",
INIT_0C => X"02E0100000000800000620100000000800000001C07261841840310240F070C3",
INIT_0D => X"0680100000000800000760100000000800000435100040000000000000080000",
INIT_0E => X"00000004000000D8008000000000000001000000155000080000000000040000",
INIT_0F => X"000100EC00004002214000008000000000000200000000000094100040000000",
INIT_10 => X"000200010C000200000000000040080005800008000001000368000040000040",
INIT_11 => X"000000004008000448000040000000000001007C000008000008001D00001000",
INIT_12 => X"000000800000000001000008000017000100000000000010200002C800000800",
INIT_13 => X"0000549000027200800E271E00288400800208004804C0080000000052800800",
INIT_14 => X"454000924280D144B14041340A880EC51160525C0022510006BE1002C6150F5E",
INIT_15 => X"010C1010C1010C3010C14086980861AD447F2201D899BA403593514B59A30088",
INIT_16 => X"010448002098694C15204369E00116203445E3443043410C5010C3010C1010C3",
INIT_17 => X"180000006018000000200804010020080400002018040000600800010064E000",
INIT_18 => X"8060000001000008060180201000000040180001006008000100201804000020",
INIT_19 => X"934D964C32698000401802008060000401000008060080201004000000080201",
INIT_1A => X"0991A185145019A28A289830C700FC0A0002870BB5ED0B34504048828464B261",
INIT_1B => X"351A8D46AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8A28A28A28A28AF4C",
INIT_1C => X"8341A0D068341A0D068341A0D068341A0D068341A0D068341A0D46A351A8D46A",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8EE3EC1A0D06",
INIT_1E => X"40155080000155FF843FFEFAA84001FF5D043FEAA5D55420AA002A8000000000",
INIT_1F => X"A80010FFAE975FFAA80001EFA2AAAAA10F7D57FEAA557BE8B45A2D5555EFAAD1",
INIT_20 => X"AAAAA105555421EFFFD568AAA002EBFEBA555542000AA80001555D04174AA002",
INIT_21 => X"280021EFA2FFE8B45F78400145FF842AAAAA2AA800BA5D51555EF002AA8BFFAA",
INIT_22 => X"00003DFEF080428B455D002AABA5D2AAAAAA5D2E82000AAD568AAA557BC0155A",
INIT_23 => X"FAAAAA8BEF552E820000851554AAFFAA801FF087BC01FF5D7FEAA105D0428B45",
INIT_24 => X"FF5D0400010AA842AAAAFFD542000FFD57DF55A280154BAA2FBE8AAAF7AA821E",
INIT_25 => X"092142E00000000000000000000000000000000000000000000015410AAD17DF",
INIT_26 => X"AB6DBEDF575FFAADE02155080E85145E3803FFEFA284051D755003DE92415F42",
INIT_27 => X"851455D0A124BA002080010FFA4955C7BE8E021C71C0A28A38EBD57DE824975E",
INIT_28 => X"B505D71424AABD7F68E2FA38555F451D7EBD16FAAA002ABFEAA555F42000E2AA",
INIT_29 => X"D56DA824975C217DAA84021FFAAF5EAB55EBAE82145F7802AABAA2A480092415",
INIT_2A => X"575EFA00012ABFB6D080A3AFEF080A2FB45490E2AA824924AAA92550A07038BE",
INIT_2B => X"AAFFEAA00F7AE821D7B6A02FBC71D0E10010005F55482E3AA801FF1471C01EF5",
INIT_2C => X"0000010400BED57FFD7410E05038BE8E2DABAFFDB6FA12ABAEBDF7DAA80104BA",
INIT_2D => X"4555043FE10087BC2000552C8000000000000000000000000000000000000000",
INIT_2E => X"ABAAAD57DE1000516ABFFFFFBD75FFAAFFC0145002897555A2803FFFFAA84175",
INIT_2F => X"DEAA557BC0010AAA895555042E820BA080400010FF8017545F7AE821455D2CAA",
INIT_30 => X"2AAAAAA8002010007FC0155D5022A955FFACBFEBA5D7BD5545A2D57DEAA002EB",
INIT_31 => X"43CAB0552C97CAAFFD57DE000057C21FFAA80001FFAAD57EB55A2A880155F780",
INIT_32 => X"AA801FF5555421EF58517EAB00028A9BEF002EAABEF002EBDF45542AAAA00080",
INIT_33 => X"A90FDFEFA280020BAA2FFEAA10FFAE82145F7803CFE55D2CC2000087BD5410AA",
INIT_34 => X"000000000000000000000002000FFD57DF55082E974AAFFAABDEBAF7FDDE6A0A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000080000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A337A20E07C0C1E006",
INIT_01 => X"295FBC448000804C5C6A60000C34C26841280A00084000C8C212802EE2953235",
INIT_02 => X"C809AD5EB118E640A4D158FC011FF0002080000082E8C66609DB7DDDCB1FA036",
INIT_03 => X"4A120E4C3A4C90D214A35E824852857A0A20640A88800000B8E0FC52A884500E",
INIT_04 => X"001440809A2604005934800041110A71E290E8B010DB221C662AE22DC0AA3448",
INIT_05 => X"12026A2A1B88C31841CDC451B860A6507BEBD18A65AE10571450DE8112522449",
INIT_06 => X"80752C03736281D628398CD0A4C894EA2054237F271331095100D82D0C2C82A2",
INIT_07 => X"5E64B66BD6231CC81529A356AD3AC601C57FF54FF149A46490261C4B39203F70",
INIT_08 => X"AD0099410015814FC602C4B1B93947F8621030C800001D7FA46A95172E937835",
INIT_09 => X"2C836D35B68D26C082DE9AB88C104020000208401807B78739010C04E17F5014",
INIT_0A => X"082099129008F25615C3FC01A2102109204C28B6706168128920C469E7C00A00",
INIT_0B => X"E92C23E210A0B246C2234010A108D0042811461C0401502644A40106C14FD22A",
INIT_0C => X"E00BF1BFE1F000BE1FC40BF1BFE1F000BE1FC80028120800800100653FF0313F",
INIT_0D => X"040BF53FE1F000BE1FC40BF53FE1F000BE1FCC806FFFEF0AE83080E2AEF2F1F1",
INIT_0E => X"013879FAAF8FC003FEDF5F12F0380231F0FF963F00A7FBDF3669C0E008C3CBFF",
INIT_0F => X"F2008022CBAC8B9DDEB779BEA91F30180309A0F83FEAB8FC7C006FFFDF1A7806",
INIT_10 => X"4131BF940DFFFE03F00003F03FB929E9C19BE8EB0C2098DFE2EF7B2760483137",
INIT_11 => X"3080E29F3B69E9F4427EEED41C0E004C72FEC95DEFE46C090626FF1537F15618",
INIT_12 => X"FC0E0392A0024B83F07F7989E9F01DFFFB0A3C0202B877EAA7A7C1CBFFD07870",
INIT_13 => X"C0404020040001C4E7F1787E0C8028514885C566241902508C83A7D1B7EFAC6D",
INIT_14 => X"4DF46A170F92C7E20F0430938008AC38C4184B100136858C9298A8560688F4C1",
INIT_15 => X"6B8C86B8CE6B8CA6B8CC15C6435C670C10EB4124D2B3903BF5C9710C1191DCA0",
INIT_16 => X"2030461200984D041C40208400230E71B3104E5636E3178C86B8CC6B8CA6B8CE",
INIT_17 => X"0040118401184610042110401184410846110421104010844118421504238200",
INIT_18 => X"8441184011844100461004211046100461084211042100441084011842100461",
INIT_19 => X"DA6924965B4D1004610840118401084410840110421004610046110421084410",
INIT_1A => X"FF9FBFAF2DDA3B9E79E7BED9CFEF73B6FFE74FC3F78FFF6DB7ED438A183124B2",
INIT_1B => X"DDEEF77BBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEDFD",
INIT_1C => X"BDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BB",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF853FB5EEF77B",
INIT_1E => X"020AA002AAAABA555140155087FFFFEF00042AB555D2E955FFF7FFC000000000",
INIT_1F => X"E975FF5D5568B555D7BD5545FFD540155FF843FFEFAA84001FF5D043FEAA5D04",
INIT_20 => X"FFEAA10F7D57FEAA557BE8B45A2D5555EFAAD5401550800001FF5D00001555D2",
INIT_21 => X"FAE975FFAA80001EF002AAAABAF7D168A10A2D17FF45A2FFC0000AAAE974AAFF",
INIT_22 => X"F7803DF55FFAEBFE005D2EAAB45557BD55555555401555D04174AA002A80010F",
INIT_23 => X"5552E955EF5D7FEAA105555421EFFFD568AAA002EBFEBA555542000A28028BFF",
INIT_24 => X"AAA2AA800BA5D51555EF002AA8BFFAAAA820AA5D517DF55082E974BA087FE8B5",
INIT_25 => X"5C7F7FBC0000000000000000000000000000000000000000000000145FF842AA",
INIT_26 => X"51D755003DE92410F42092142E28ABA5D5B4516D007FFFFFF1C042FB7D492A95",
INIT_27 => X"851C75D0E02145492E955C75D5F6DB55497BD5545E3DB45145E3803AFEFA2840",
INIT_28 => X"BC7028A2AA95492FFFFE8A38EBD57DE824975EAB6DBEDF575FFAADF42155082E",
INIT_29 => X"0A124BA002080010FFA4955C7BE8E021C71C0A2DABAF7D16DA28A2DB7AF7DB6F",
INIT_2A => X"55F42000E2AAA8BEFE3843AF55E3AABFE105520AFB45557BD5555415F4514549",
INIT_2B => X"082E954AA087FEDB7D5D2A155D7157BEFA38555F451D7EBD16FAAA002ABFEAA5",
INIT_2C => X"0000002145F7802AABAA2A480092415B505D71424821D7F68E07082495B7FF7D",
INIT_2D => X"EF5D003DFEF002E95555F7FDC000000000000000000000000000000000000000",
INIT_2E => X"555A2802ABFFAA841754555043FE10082A82000552CAAAAA5D7FD75EF087BFDF",
INIT_2F => X"75FFAAFFC0145002895545552E80145002E955455D7BFDF45007FD7555A2F9D5",
INIT_30 => X"7FEAAAAFFEABFFF7FFD54BAA2AA95410F7FDEAABAAAD57DE1000516ABFFFFFBD",
INIT_31 => X"BD55550879D5555002E820BA080400010FF8017545F7AE821455D2CBFEAAFFD1",
INIT_32 => X"D57DEAA002EBDEAA557BC0000AAA8A8BEFA28028B45AAAABFE0009043FF555D7",
INIT_33 => X"FAC97400087FFFFFF002E954AA087BFFFFF5D2E975455D7DFFEBA5D7BD5545A2",
INIT_34 => X"000000000000000000000000155F7802AAAAAA8002010007FC0155550222955F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000300000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B0061A258A2840112C03002C180004003220200403302301C0381A0082",
INIT_01 => X"860041C838394848008100000042026041000000090800090210010000510204",
INIT_02 => X"080108220C1000004464080000C008010000000001243240080080000988A050",
INIT_03 => X"080000010C23404080020A600200002983800504488000103080050C08C10000",
INIT_04 => X"0040504280A682104011230010000010002040E9102050101000400A00003000",
INIT_05 => X"0409400984008000414A00014000002004100020005004020010204044802800",
INIT_06 => X"301223FC028911E8911900000224200248A653E908C0248489FF000809108000",
INIT_07 => X"0000220441820000090C080001184400142040200E824008900008000220600A",
INIT_08 => X"1A18946451007FA0380200808809010C182000000000090F8100001220000804",
INIT_09 => X"300240B4A409223F020988100808200490142B441BF82C20401481540A000008",
INIT_0A => X"264285180542408000D001BE090693912000002004410489080001100017E2FD",
INIT_0B => X"091081090A4491A40052A129519428CA142288010A5A21214601F01A220602A0",
INIT_0C => X"18100400000000A00034100400000000A00033A00813004104020818800F2400",
INIT_0D => X"F4100080000000A00034100080000000A0003142000000000000000000055D00",
INIT_0E => X"00000001E8002900010000000000000000066000C20004000000000000000120",
INIT_0F => X"4D240C2000502000000080000000000000000000240146800142000000000000",
INIT_10 => X"00001260F0000000000000000007F00032201000000000091A00040000000002",
INIT_11 => X"0000000005D00008958010000000000000003F4000008000000048D240008000",
INIT_12 => X"008000000000000000082670000CC0000000000000000007C000301400200000",
INIT_13 => X"0120849A5250101482202301F05101202420000810C219500150002800101280",
INIT_14 => X"454110030212C140011204D020880C000018431DE802015022A62A1596C8B580",
INIT_15 => X"016C2016C2016C6016C440B6000B600C446B0104D09192013589701C59800002",
INIT_16 => X"51804A0028904C425016040820978221B0000005B05B416C0016C0016C4016C4",
INIT_17 => X"8CA3294A528CA328CA1294A528CA3284A5294A728CA3284A529CA728CA100508",
INIT_18 => X"CA3284A129CA7294A328CA1294A729CA128CA329CA5294A128CA3294A5294A32",
INIT_19 => X"1C71C718638E28CA529CA7284A128CA7294A528CA1284A729CA1284A3284A529",
INIT_1A => X"ED9DBDAFBC5E9BBEFBEFBEF9CFF1FE1E9F52AFF9F3E77B7CF7F40A00107638C3",
INIT_1B => X"FCFE7F3F8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E76C",
INIT_1C => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9",
INIT_1D => X"00000000000000000000000000000000000303007FFFFFFFFFFFC61AC8FE7F3F",
INIT_1E => X"955FFF7FFC21EFF7D17DEAA5D2AAAAAA5D557DE105D2EBDF55557FC000000000",
INIT_1F => X"03DEAA5D5568BEF5D042AA10A2AAAAABA555140155087FFFFEF00042AB555D2E",
INIT_20 => X"5540155FF843FFEFAA84001FF5D043FEAA5D00020AA002A82145555542010FF8",
INIT_21 => X"D5568B555D7BD5545FFD568AAA5D00154AAAAD1420BA00557DF455D7BFFEAA55",
INIT_22 => X"F7843FF55007FFDEAAA284020BAAAD168BFF0800001FF5D00001555D2E975FF5",
INIT_23 => X"5AAAEBFE10FFFFEAA10F7D57FEAA557BE8B45A2D5555EFAAD540155080000000",
INIT_24 => X"10A2D17FF45A2FFC0000AAAE974AAFFFFC21EF5551401EFF7842AA00FF841754",
INIT_25 => X"F45497FC000000000000000000000000000000000000000000002AABAF7D168A",
INIT_26 => X"FFFF1C042FB7D492A955C7F7FBC71EFFFD57FE825520ADA92495B7AE10412EBF",
INIT_27 => X"0716D415F47000F78A3DE92415F6ABD7490A28A10AAAAA8ABA5D5B4516D007FF",
INIT_28 => X"F78F7D497FFFE925D5B45145E3803AFEFA284051D755003DE92410E02092140E",
INIT_29 => X"0E02145492E955C75D5F6DB55497BD5545E3DB6AA92550A104AABED1470AA005",
INIT_2A => X"ADF42155082E87038FF8038F6D1C7BF8EAAAA80020BAA2DB68BC7140E051C75D",
INIT_2B => X"FF8428A00E38412545AAAE3FE10A3FBE8A38EBD57DE824975EAB6DBEDF575FFA",
INIT_2C => X"000002DABAF7D16DA28A2DB7AF7DB6FBC7028A2AA95492FFFFC71EF415F471C7",
INIT_2D => X"00007FEAA10002ABFF450079C000000000000000000000000000000000000000",
INIT_2E => X"AAA5D7FD75EF087BFDFEF5D003DFEF002E95555F7FDD55EFF7D57DE005D003DE",
INIT_2F => X"FE10082A82000552C955FF007BD5410FFAABFE00087BE8B45082EAAA10A2A8AA",
INIT_30 => X"820AAF7D5574AA087BEABEF007FFDE00557DD5555A2802ABFFAA841754555043",
INIT_31 => X"BEAB55552C95545552E80145002E955455D7BFDF45007FD7555A2F9EAA005D2A",
INIT_32 => X"516ABFFFFFBD75FFAAFFC01450028974BAFF842ABFF557BE8ABAA284020BAA2F",
INIT_33 => X"7FDD55EF007BD5555F7802AA10AA8000145AAAEBFE10A2F9EAABAAAD57DE1000",
INIT_34 => X"00000000000000000000003FEAAFFD17FEAAAAFFEABFFF7FFD54BAA2AA95410F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000240000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C024504188000003000000003302300C018180006",
INIT_01 => X"020008422008604D042080000211024840000000080000080200080000110204",
INIT_02 => X"4801082048100000444008040080000041000000000222400800000009000010",
INIT_03 => X"0802030288A148D0000208424000002103006400088000003080000408C10000",
INIT_04 => X"00004000890600004032030010000010008060E4100000140006500800403040",
INIT_05 => X"0400400080000018414800810000002000000000004000328010000080882000",
INIT_06 => X"281A8001220021E0021803000224200200000360888420000000100808000000",
INIT_07 => X"5000220409020000090800000118040014A061200052500810000C490323208E",
INIT_08 => X"1A9098411110014000424090980B0002102000000000010F8000001220000805",
INIT_09 => X"31024034A4092200820D899408000004D0143B4410002C800080020450800001",
INIT_0A => X"24028011444240A88CC00100200D0010200008B2066397014800221400140C01",
INIT_0B => X"080001000C008124000000000100008000100404204C25200451A01A00A620A5",
INIT_0C => X"1C0014800000F001E02C0014800000F001E021141213000000000010B0001000",
INIT_0D => X"CC0014800000F001E02C0014800000F001E022420000400004C3201C51040908",
INIT_0E => X"60078601084038000180400002C0E00E0E004100E000040900000B0380383400",
INIT_0F => X"08146800105100000000800284004160C0301D07001504820242000040000198",
INIT_10 => X"908C404AFC000200030F000FC00610103BE0104810C8462014F8040446120C88",
INIT_11 => X"C3201C608410100FD5801044013098038D00309F008088C2419100A7C0209021",
INIT_12 => X"00B2048902C0807C0E008450100FDD000100411C8107880440403DDC00201804",
INIT_13 => X"00100496406010A0A2002200125140000000221110C018066250402E32901A80",
INIT_14 => X"454214028220141530400910CA800900326790500002001444001C0050140A00",
INIT_15 => X"5120551205512055120708901A8901A104804000801212541403C15178008010",
INIT_16 => X"01004200A09A49445420000DC000152804C9A384814809201512015120151201",
INIT_17 => X"0004000000080200806008020000000000000020080200802000000000008000",
INIT_18 => X"0000000000802008000000000002008020000400000000000080600802008000",
INIT_19 => X"0002082080000100000802008020100000000008020180000000000020180200",
INIT_1A => X"0000000000000000000000000000000000000000000000000005428A14584104",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8DD9EC000000",
INIT_1E => X"BDF55557FFDE00557BEAABAA2AEAABEFF78015555AA801741055554000000000",
INIT_1F => X"BEAAAAAAD157555AA803FEBA5555421EFF7D17DEAA5D2AAAAAA5D557DE105D2E",
INIT_20 => X"802AABA555140155087FFFFEF00042AB555D2E955FFF7FFD5555557BEABFFF7F",
INIT_21 => X"D5568BEF5D042AA10A2AA955EFF7FFD5400F7FFFDFEFAA80000BAAAAA820BAA2",
INIT_22 => X"5D7FE8A000004154BAF780001EFAAAAA8B45000002145555542010FF803DEAA5",
INIT_23 => X"5AAD5555EF557FC0155FF843FFEFAA84001FF5D043FEAA5D00020AA002ABDEBA",
INIT_24 => X"AAAAD1420BA00557DF455D7BFFEAA5555575455D2AAABFF5551421FFAAD15754",
INIT_25 => X"4385D5540000000000000000000000000000000000000000000028AAA5D00154",
INIT_26 => X"DA92495B7AE10412EBFF45497FFFE385D71E8AAAAAA0A8BC7EB8417555AA8410",
INIT_27 => X"D056D5D75EABC7FFF5EAAAABEDF5257DAA8438EBA4155471EFFFD57FE825520A",
INIT_28 => X"0070BAA2A0870BAAA8028ABA5D5B4516D007FFFFFF1C042FB7D492A955C7F7FB",
INIT_29 => X"5F47000F78A3DE92415F6ABD7490A28A10AAAA925EFEBFFD2400EBFBFAFEFAA8",
INIT_2A => X"10E02092140E3DE924171E8A281C0E10482F784001D7AAA0AFB6D1C040716D41",
INIT_2B => X"4955421EFA2DF5557DAAD5D05EF0175C5145E3803AFEFA284051D755003DE924",
INIT_2C => X"000002AA92550A104AABED1470AA005F78F7D497FFFE925D5B525454124AFBC7",
INIT_2D => X"55A28015545A284000BA5D534000000000000000000000000000000000000000",
INIT_2E => X"5EFF7D57DE005D003DE00007FEAA10002ABFF450079FFEAA5D5568ABAA2842AB",
INIT_2F => X"DFEF002E95555F7FDC01EF55556AB55F7D56AABAF7FBC01EFA2842AABA085755",
INIT_30 => X"C2000A2FFEABFFAA84174BAAA80174AAAA862AAAA5D7FD75EF087BFDFEF5D003",
INIT_31 => X"43DFEF5D02155FF007BD5410FFAABFE00087BE8B45082EAAA10A2A8801FFA2FF",
INIT_32 => X"841754555043FE10082A82000552CBFE10085168AAA552A80010F78000145AA8",
INIT_33 => X"57DC014500003FF450051401FFA2FBD55EFAAD5421FF085755555A2802ABFFAA",
INIT_34 => X"00000000000000000000002AA005D2A820AAF7D5574AA087BEABEF007FFDE005",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0000040042840002C00000018000002700500030B3132000400812082",
INIT_01 => X"A14008420008204D042100000212026840000000180800080200090048510200",
INIT_02 => X"080108020090000004655C000080000051000000002402400800000009008010",
INIT_03 => X"0002000100300C408422420002108108028065044880001030808D4288C10000",
INIT_04 => X"0002504688A28210003100000000001002A0E88910A032541000090A00643040",
INIT_05 => X"04092A081400D118410A002140004020140001A9005000004810A1C0044D2800",
INIT_06 => X"0010EFFD228931C8931820002080258A48A653E00213248C98FFC0094910A222",
INIT_07 => X"4000220440120000090C0810210A040034A040000046180810000C4907036008",
INIT_08 => X"50D88C2450000140004200808809000C012000000000010F8102041320000000",
INIT_09 => X"2002002020010200828C88020800200040801A40100228A1585481544A804040",
INIT_0A => X"A20804802400C80080D0010029069290200008B20E2304086800400640200801",
INIT_0B => X"091084090A4C81240251A328D094684B34A288050A5828012009504420102180",
INIT_0C => X"080004801E0FF00010000004801E0FF000100220021200000000000080001000",
INIT_0D => X"000004801E0FF00010000004801E0FF000100440000000F517CF600000400104",
INIT_0E => X"E000004008100800010040ED0FC7E000004008804000040109963F1F80000080",
INIT_0F => X"0020040020100000000882431660CFE7C0F00000000800810040000000E587F9",
INIT_10 => X"B0000808000001F80FFF0000200008021040134473D800040010045C1F360001",
INIT_11 => X"CF600000200802028001102EA3F1F80000400002008B83D6C0002000802688E7",
INIT_12 => X"03F2DC2D1FC18000000040080202800004D5C3FD80000080200818000027928F",
INIT_13 => X"0122C01A52501094222002000110012064200008848218002100100C00004112",
INIT_14 => X"4500048240C08400841204D0A00089000100001DE9248104300294428148A480",
INIT_15 => X"4800048000480004800004002240020850884000901210140011C010312B888A",
INIT_16 => X"51A4C000889A4D0E1D7624086491800420044240020004004480004800048000",
INIT_17 => X"84A1284A128CA328CA328CA328CA328CA328CA1284A1284A1284A12C4A14E508",
INIT_18 => X"CA328CA3284A1284A1284A1284A328CA328CA328CA328CA3284A1284A1284A12",
INIT_19 => X"000000000000284A128CA328CA328CA328CA3284A1284A1284A1284A328CA328",
INIT_1A => X"4799B1A014503EB65B6594F14A87D78AF421448BB528AF75D640088884400000",
INIT_1B => X"7C3E1F0F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79EDFC",
INIT_1C => X"87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F0F87C3E1F0F8",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF834FA53E1F4F",
INIT_1E => X"174105555420000000021EFAA843DE00F7803FEBAFFFFC2000557FC000000000",
INIT_1F => X"43DE005504175FF08514014555557DE00557BEAABAA2AEAABEFF78015555AA80",
INIT_20 => X"7FC21EFF7D17DEAA5D2AAAAAA5D557DE105D2EBDF55557FD54AAA2AA955FF000",
INIT_21 => X"AD157555AA803FEBA55556ABFFA280154BAFF803DF45FFD17DFFFFFD56AA0055",
INIT_22 => X"002AAAAAAA2D57DF450004154BA087BEAAAAF7D555555557BEABFFF7FBEAAAAA",
INIT_23 => X"5FFD1555EFA2802AABA555140155087FFFFEF00042AB555D2E955FFF7FFD5410",
INIT_24 => X"00F7FFFDFEFAA80000BAAAAA820BAA280000AAA2843DE1008556AA00A28028B5",
INIT_25 => X"0285D75C00000000000000000000000000000000000000000000155EFF7FFD54",
INIT_26 => X"8BC7EB8417555AA84104385D5542038000A001C7A2803AE38FF843DEBAEBFFC2",
INIT_27 => X"D24BAA2AA955C708003FE285D00155FF0055451555D5F7FE385D71E8AAAAAA0A",
INIT_28 => X"B78FFFE3DF6DA284175C71EFFFD57FE825520ADA92495B7AE10412EBFF45497F",
INIT_29 => X"75EABC7FFF5EAAAABEDF5257DAA8438EBA415568BEFA28E124AAF7843AF7DEBD",
INIT_2A => X"92A955C7F7FBD54380020ADA82BED57DF450804104920875EAA82F7DB5056D5D",
INIT_2B => X"005F68A10BE802DB55E3DB555FFF68028ABA5D5B4516D007FFFFFF1C042FB7D4",
INIT_2C => X"00000125EFEBFFD2400EBFBFAFEFAA80070BAA2A0870BAAA80070BAA2803DE00",
INIT_2D => X"AAFF803DEBAAAFBC20BA55514000000000000000000000000000000000000000",
INIT_2E => X"EAA5D5568ABAA2842AB55A28015545A284000BA5D53420BA082E82155AA802AA",
INIT_2F => X"AA10002ABFF450079C20BAAAAE9754500043DEBA5D04175EF0855575455D7BFF",
INIT_30 => X"820AAFF802ABEFAAFFEABEFAAFFFDEAA0051555EFF7D57DE005D003DE00007FE",
INIT_31 => X"16AA10FFFFC01EF55556AB55F7D56AABAF7FBC01EFA2842AABA085768BFFA2AE",
INIT_32 => X"7BFDFEF5D003DFEF002E95555F7FDD74BA08043DE10F7D17FF55000000010085",
INIT_33 => X"A86174AAAA843DE00087FE8A00F7843FF45AAFFD75EFF7842AAAA5D7FD75EF08",
INIT_34 => X"0000000000000000000000001FFA2FFC2000A2FFEABFFAA84174BAAA80174AAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000100000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000006",
INIT_01 => X"000009801830084C182060000C104268413C0A61590001D90213C00000110200",
INIT_02 => X"680108200010000054400C000080000041000000010002400800800009082011",
INIT_03 => X"0008000004002040000200100000000042800584488000103081880008800000",
INIT_04 => X"00005842802AC210001000000800001000004080100040140080040800003100",
INIT_05 => X"0400000040000080410800010001002000000000004000002010000040002000",
INIT_06 => X"10100001221911E1911902000020200201A2D3E8000C2C84880010080800004C",
INIT_07 => X"C0002204000200000B080000010C040004A0400000C0000810000C5901036000",
INIT_08 => X"002A84300000014000C2008088090000002000000000030F8000001220000408",
INIT_09 => X"210000020000120082088801080020400000084010002880000C803400000008",
INIT_0A => X"020000040000480100D0010019019190200008B2022380800802010000000801",
INIT_0B => X"09000119064C810500D0A36851B428DA14368C801A1400000100500400000090",
INIT_0C => X"08100080000000A00000100080000000A00000000212000000000000B0001000",
INIT_0D => X"00100400000000A00000100400000000A0000540000000000000000000005100",
INIT_0E => X"00000000A8000900000040000000000000060000420000010000000000000120",
INIT_0F => X"4000040000102000000000020000000000000000240000800140000000000000",
INIT_10 => X"00001204FC000000000000000001280013A000400000000900E8000400000002",
INIT_11 => X"0000000001480004D5800004000000000000091D008000000000480740200000",
INIT_12 => X"0002000000000000000820080004DD000000000000000002A00011DC00001000",
INIT_13 => X"0322C01032301006022082000010032024200000048019500000000832901A80",
INIT_14 => X"4501000200089400007200D0020008000000144C4800000200BC228404020080",
INIT_15 => X"0010000104001000010440080000822900000000801010500A13404111008000",
INIT_16 => X"D1A0CA0000984D06403600086591900224002000400440104001040010000104",
INIT_17 => X"8DA368DA3685A1685A1685A1685A1685A1685A1685A1685A1685A1685A120D08",
INIT_18 => X"5A1685A1685A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA36",
INIT_19 => X"000000000000685A168DA368DA368DA368DA368DA368DA368DA368DA1685A168",
INIT_1A => X"6C20080AB9A28724904120E1999E91BCD151200802001038E2550A0010100000",
INIT_1B => X"68341A0D14514514514514514514514514514514514514534D34D34D34D344A1",
INIT_1C => X"268341A0D069349A0D069349A0D068341A4D268341A4D268341A0D068341A0D0",
INIT_1D => X"00000000000000000000000000000000000003FFFFFFFFFFFFFF8A6AC8341A4D",
INIT_1E => X"C2000557FEABEFA2D1400AA5D2AAAA00F7FFEAA10F7D17FFFFAAAE8000000000",
INIT_1F => X"03DFEFF7FFE8ABAF7802ABEFAAAE820000000021EFAA843DE00F7803FEBAFFFF",
INIT_20 => X"843DE00557BEAABAA2AEAABEFF78015555AA80174105555421EFF78028BEF5D0",
INIT_21 => X"504175FF0851401455555555EFA2FBC01FFF7AAAAB45557BC0155007FFDEBAAA",
INIT_22 => X"552A974AAA2843DEAA5D2A820BA000428AAAAA84154AAA2AA955FF00043DE005",
INIT_23 => X"AF7D1400BAAAAE821EFF7D17DEAA5D2AAAAAA5D557DE105D2EBDF55557FFDE00",
INIT_24 => X"BAFF803DF45FFD17DFFFFFD56AA00557FC201000517FFEFAAAEBDF45FFAEA8AB",
INIT_25 => X"FD7A2A48000000000000000000000000000000000000000000002ABFFA280154",
INIT_26 => X"AE38FF843DEBAEBFFC20285D75EFBC7A2DB400824120ADA38E3F1EFA28F7DF7D",
INIT_27 => X"421C7FF8028BEF41003FFD7F7F1EDA82F78E2DBD7A2A482038000A001C7A2803",
INIT_28 => X"1C716D1475FFEAAA28E3FE385D71E8AAAAAA0A8BC7EB8417555AA84104385D55",
INIT_29 => X"AA955C708003FE285D00155FF0055451555D5F575C7A2FBC51EFEBA0A8B6D557",
INIT_2A => X"12EBFF45497FFFE105D2E97482AA8038EAA412E850AA1C0428ABAB68E124BAA2",
INIT_2B => X"B6A0BFF55F7AEAAA82FFDF40092B6A4871EFFFD57FE825520ADA92495B7AE104",
INIT_2C => X"0000028BEFA28E124AAF7843AF7DEBDB78FFFE3DF6DA284175C001000557FFEF",
INIT_2D => X"AAA2D57FEAAF7FBFDF45AA800000000000000000000000000000000000000000",
INIT_2E => X"0BA082E82155AA802AAAAFF803DEBAAAFBC20BA55517DF55A2FBC201008003DE",
INIT_2F => X"5545A284000BA5D5340145F78028BFF08003DF45FFD57FE00FFAABFF45AA8002",
INIT_30 => X"D75FFA2842ABFF5555575FF55557FEAAA2AABFEAA5D5568ABAA2842AB55A2801",
INIT_31 => X"028ABAF7AA820BAAAAE9754500043DEBA5D04175EF0855575455D7BD5555A2FB",
INIT_32 => X"003DE00007FEAA10002ABFF450079FFE005D2A97400A2802AABA002A954AA5D0",
INIT_33 => X"0514200008517DFEFFF803FF45FFAAA8A00F7FBC2010FF80155EFF7D57DE005D",
INIT_34 => X"000000000000000000000028BFFA2AE820AAFF802ABEFAAFFEABEFAAFFFDEAA0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000200000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110204",
INIT_02 => X"0801080200100000046558040080000041000000002402400800000009008010",
INIT_03 => X"00020201040000D0842242024210810802006400088000003080054288C10000",
INIT_04 => X"0000400088020000003020002000001002A0E881108032100002000800203040",
INIT_05 => X"04092A081000411841480001000000201000012800400010001081C040402000",
INIT_06 => X"10100001220001E0001802002020240208000369001520080100100909000266",
INIT_07 => X"4000220440020000090C0810210A040004A0410000C0000810000C4901036008",
INIT_08 => X"0000802100100140004200808809000C002000000000010F8102041320000000",
INIT_09 => X"2000000000000200828888800808000410800840100220211850004442004048",
INIT_0A => X"240A80800442400004C0010000060210200008B2022304880800410000200801",
INIT_0B => X"0000010008008020020100008000400120800004004821202001A05A00040180",
INIT_0C => X"08101400000000A01004101400000000A0100000081300410402080080003000",
INIT_0D => X"04101080000000A01004101080000000A0100540000040000000000000405100",
INIT_0E => X"00000040A80009000180000000000000004608004200040800000000000001A0",
INIT_0F => X"4000282000102000000080008000000000000000240800800140000040000000",
INIT_10 => X"00001A00000002000000000020013000100010080000000D0000040040000003",
INIT_11 => X"0000000021500000800010400000000000400900000088000000680000009000",
INIT_12 => X"008000800000000000086010000080000100000000000082C000100000200800",
INIT_13 => X"040004924040008020000200101100004000000000C019500050000800000000",
INIT_14 => X"4541008240801000804000108280800001001051A12481041080801010000080",
INIT_15 => X"4800048004480044800044000240022100884000901210440003C141102B088A",
INIT_16 => X"00044280009048485D4020080000140004046240020044000480044800448000",
INIT_17 => X"080200802008020080200802008020080200802008020080200802048026E011",
INIT_18 => X"0000000000000000000000000002008020080200802008020080200802008020",
INIT_19 => X"0000000000000080200000000000000000000000000000000000000000000000",
INIT_1A => X"CA83332A34488A8A28A29E195281FC1A72E24C2BF5A4D9555204428290100000",
INIT_1B => X"94CA65328A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A354",
INIT_1C => X"994CA6532995CAE572B94CA6532994CA6572B95CAE532994CA6532994CA65329",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF838CF1CAE532",
INIT_1E => X"7FFFFAAAE801FF08557DF4555516AA00007BEABEFAAD1555FFF7840000000000",
INIT_1F => X"56AA0000043FFEFA2FFFDE1008556ABEFA2D1400AA5D2AAAA00F7FFEAA10F7D1",
INIT_20 => X"84020000000021EFAA843DE00F7803FEBAFFFFC2000557FC0010AAD57FF45A2D",
INIT_21 => X"7FFE8ABAF7802ABEFAAAEA8BFF5D0415400F7FBFDEAA007FEAB45AAAE800AAF7",
INIT_22 => X"5D0415555557BFDFEF00517DE00A28028B450855421EFF78028BEF5D003DFEFF",
INIT_23 => X"A5D7FFDEBAF7AEBDE00557BEAABAA2AEAABEFF78015555AA80174105555401FF",
INIT_24 => X"FFF7AAAAB45557BC0155007FFDEBAAA8417410AAFFD7555AAD56AB45A2AE800A",
INIT_25 => X"5C7E380000000000000000000000000000000000000000000000155EFA2FBC01",
INIT_26 => X"DA38E3F1EFA28F7DF7DFD7A2A4801EF085F7AF6D55556AA381C75EABEFBED157",
INIT_27 => X"C0010AADF7AF6DB6D56FA3814003AFFFA2F1F8E381C516FBC7A2DB400824120A",
INIT_28 => X"5E8B45BEA0850BAE38002038000A001C7A2803AE38FF843DEBAEBFFC20285D75",
INIT_29 => X"8028BEF41003FFD7F7F1EDA82F78E2DBD7A2A4ADBEF550412428F7F5FDE92087",
INIT_2A => X"A84104385D55401C75504125455575FAFD7145578E10AA802FB450851421C7FF",
INIT_2B => X"BED56FB45BEA082082557BF8EBAF7AABFE385D71E8AAAAAA0A8BC7EB8417555A",
INIT_2C => X"00000175C7A2FBC51EFEBA0A8B6D5571C716D1475FFEAAA28E10438AAF5D2545",
INIT_2D => X"BA5D5568BEFF7D157555AA800000000000000000000000000000000000000000",
INIT_2E => X"F55A2FBC201008003DEAAA2D57FEAAF7FBFDF45AA80021FF007BE8BFF5D516AA",
INIT_2F => X"DEBAAAFBC20BA555140010AAFFE8BFFFFD17DEBA5D002ABFFA2D16AAAA55517D",
INIT_30 => X"020BAFFD17DE10005568B55FF80154BAA280020BA082E82155AA802AAAAFF803",
INIT_31 => X"43FF55085140145F78028BFF08003DF45FFD57FE00FFAABFF45AA803FFEF5500",
INIT_32 => X"842AB55A28015545A284000BA5D53421455504021555D556AB555D5568A00AA8",
INIT_33 => X"2AA800AAAAD142155F7D57DF45FF8002010557FEAAAAF7AABFEAA5D5568ABAA2",
INIT_34 => X"000000000000000000000015555A2FBD75FFA2842ABFF5555575FF55557FEAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000023FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B83008481800E0000C26426040000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"00080D4912E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"000048048002400048150000000002504230C899109032100020160880223000",
INIT_05 => X"040B2A229100410041088011100022201200012840440000B01088C0005C2400",
INIT_06 => X"287E4003225021C5021880C02000A40249048363A5992808110010090908022A",
INIT_07 => X"4044222987020C80152D8910210A0400252B74200045C86810000C5B0503286A",
INIT_08 => X"26509804400501400242C0B0B83B0134702000000000191FA162841324832069",
INIT_09 => X"3002000220001240820F8B2A08000040409018401001200159D80D64AA004041",
INIT_0A => X"020808852000420718C00101B0070310200008B60A23A51B2802467327200801",
INIT_0B => X"080802500C08832582810240812040912094068010050402214850444091019B",
INIT_0C => X"761B011986695014A96E1A8119865A5018C5A0A00012004104020808B0003000",
INIT_0D => X"AE1A811986695014A96E1B0119865A5018C5AF0062C38A4DB680A0D8241501D5",
INIT_0E => X"802CAB184E8F4101621B1BAC845542056A289A1BB2078A922DA2A8B180A2600A",
INIT_0F => X"392000224ACDE215883078681B5C05AA429189B60AC43CEC7F0272C3841DB528",
INIT_10 => X"51BCA1C90006C0C2958502861120C003104289A668B8CAB270106338317A3D94",
INIT_11 => X"A64090B89E015AAA880E48382EB8804B020A06020C67061BC785938085134CD5",
INIT_12 => X"C6284B2D20410AB4503089C00A8280819A5539D503336D61056ABA006282806C",
INIT_13 => X"060040142020015001004A00080042004000E8089C9003066E03513E41470126",
INIT_14 => X"4536708201C000908020349320008000A1000C09A9348498B000000000000080",
INIT_15 => X"32A0C32A0C32A0832A0C19504195040040000000801010028001400010010CBA",
INIT_16 => X"8104400000904C0C0964200841010954000444D280140050C32A0832A0C32A08",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090246811",
INIT_18 => X"1004010040100401004010040102409024090240902409024090240902409024",
INIT_19 => X"0000000000004010040100401004010040100401004010040100401004010040",
INIT_1A => X"488292A831308E0000000A11100830181621409A14E871104201400284000000",
INIT_1B => X"0000000000000000000000000000000000000000000000020820820820820A05",
INIT_1C => X"0000000402000000000000000000010080000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8C0F00000000",
INIT_1E => X"555FFF784020AAF7D542155F7D1400AAF7FFFDE00F7842AA00002A8000000000",
INIT_1F => X"A800AA007FFDFFFA28428A000000001FF08557DF4555516AA00007BEABEFAAD1",
INIT_20 => X"FBEABEFA2D1400AA5D2AAAA00F7FFEAA10F7D17FFFFAAAEA8ABAFFD17FEBAFFA",
INIT_21 => X"0043FFEFA2FFFDE1008556AB45555568A10A2FFC00AAF78028AAAFF84020AAFF",
INIT_22 => X"FFD1555FF0804000AA000428A10AAAA801EFFFD140010AAD57FF45A2D56AA000",
INIT_23 => X"FA2FBFFF550000020000000021EFAA843DE00F7803FEBAFFFFC2000557FC0155",
INIT_24 => X"00F7FBFDEAA007FEAB45AAAE800AAF78428B45A28428A10087FD7400552EBDFE",
INIT_25 => X"A101C2A80000000000000000000000000000000000000000000028BFF5D04154",
INIT_26 => X"AA381C75EABEFBED1575C7E380000BAF7DB4016DE3DF450AAF7F1FDE38FF8A2D",
INIT_27 => X"AFABAFFDF7AE82F7AA870AA0071F8FFFBE842DA101C0E001EF085F7AF6D55556",
INIT_28 => X"42DAAAE38A02082E3FBEFBC7A2DB400824120ADA38E3F1EFA28F7DF7DFD7A2A4",
INIT_29 => X"DF7AF6DB6D56FA3814003AFFFA2F1F8E381C516DB455D5B68A28A2FFC20AAEB8",
INIT_2A => X"BFFC20285D75C2145F7DF525EF140A050AA1C0028A28AAA4801FFE3DF40010AA",
INIT_2B => X"007FD74284120BFFFFBEF1F8F7D080A02038000A001C7A2803AE38FF843DEBAE",
INIT_2C => X"000002DBEF550412428F7F5FDE920875E8B45BEA0850BAE3802DB6DAA8A28A00",
INIT_2D => X"AAF7D57DEAAF7AABDE10552E8000000000000000000000000000000000000000",
INIT_2E => X"1FF007BE8BFF5D516AABA5D5568BEFF7D157555AA80020BAFFFBC01EFA2FFD74",
INIT_2F => X"FEAAF7FBFDF45AA803FEBAFFFBEAA00F7AE974BA085568BEFF7803FE10552E82",
INIT_30 => X"EAAAAA2FFC00AAAA803FEAAA2AA82000A2FFFDF55A2FBC201008003DEAAA2D57",
INIT_31 => X"0001FFAAFFC0010AAFFE8BFFFFD17DEBA5D002ABFFA2D16AAAA55517DF55557F",
INIT_32 => X"802AAAAFF803DEBAAAFBC20BA555142155F7FFC01EF552E974BA550028ABAA28",
INIT_33 => X"2803FFFFA2AAAAA00007FD74BA08003DFFFFFD16ABFF082E820BA082E82155AA",
INIT_34 => X"00000000000000000000003FFEF5500020BAFFD17DE10005568B55FF80154BAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000200000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702684000000008000008820009280A553231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"421A0A0012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"02004000890200001837830011998C31C09060DC104000102002140900003548",
INIT_05 => X"0402002BC200009841090001200006200800000020480010A4100100001C2000",
INIT_06 => X"287FC003230001D0001806C0060CB0622000037085C820000000100C0C200008",
INIT_07 => X"CE64B663DFA314C803292140890C0601F472D1640051F80C10020C493F033432",
INIT_08 => X"67C081000111814004C20481A92940EA7A3020480000071F846890162E135038",
INIT_09 => X"240048108488024082488BAF08000020800629441004300421800F04F8000001",
INIT_0A => X"A0200E0BF40063FF9DC0010000180018200408B27E234913E900067F04D40C01",
INIT_0B => X"002002801000A04200000000000000000000029D204B7C0382FD0100F3F9F80F",
INIT_0C => X"7E0B348EDAC3900F6EFA0B158EDA93900F6EE230381208008001007A80001100",
INIT_0D => X"CA0B158EDAC3900F6EFA0B348EDA93900F6EE8421392C96B1237E0D8BD9628F9",
INIT_0E => X"412EDD2B47CFF812A383430C669E622DBC31D73F6006A5891533EF9500EAE64B",
INIT_0F => X"BA30E022DAD8C100CA39E8CEBE66C2B083798D341B10DE7E14400392C74CAEAD",
INIT_10 => X"71A9C5DD00B12728D5360234D62A49FAB442994B3238D4E2FB104636652E19B8",
INIT_11 => X"C800DA550C29F36A8A2554E48A6430469392526208C6CC95C33717D885329664",
INIT_12 => X"51B60585A5C28895962502E9F36A828C4999AF580395542D27CDBA0020F0FABA",
INIT_13 => X"0000001E404011F066000A000EE040000000873FB80B8A00EF03F56CC12B416A",
INIT_14 => X"4D667C06CC6816B300403C13E2000000460010400000010CE080801010000080",
INIT_15 => X"72F0C72F0872F0872F0C597863978421040800209010124ACA03414158228430",
INIT_16 => X"00104280A89A4D004000000800001D5E05182493C5BC5AF0872F0C72F0872F08",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000010000",
INIT_18 => X"8020080200802008020080200800000000000000000000000000000000000000",
INIT_19 => X"0000000000000080200802008020080200802008020080200802008020080200",
INIT_1A => X"E02000028DCA05A8A28A2048C1111026C152A2316246000CB054420210100000",
INIT_1B => X"C864321904104104104104104104104104104104104104124924924924924481",
INIT_1C => X"2C964B2592C964B2592C964B2592C964B2592C964B2592C964B2190C86432190",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800FFD64B259",
INIT_1E => X"2AA00002AAAA10FF8002155F7FFC2000080417555FFAA80155F7840000000000",
INIT_1F => X"FE8AAA080000155F7FFFDEAA0000020AAF7D542155F7D1400AAF7FFFDE00F784",
INIT_20 => X"2E801FF08557DF4555516AA00007BEABEFAAD1555FFF7842AB55080000145557",
INIT_21 => X"07FFDFFFA28428A00000028B4555043DFFFFFAE82000FF80020AAA2AAAABFF00",
INIT_22 => X"A284174AAFF8428AAAFF8415545AAFBD7545F7AAA8ABAFFD17FEBAFFAA800AA0",
INIT_23 => X"5F7FFFDEAA08556ABEFA2D1400AA5D2AAAA00F7FFEAA10F7D17FFFFAAAE80000",
INIT_24 => X"10A2FFC00AAF78028AAAFF84020AAFFFBC21550800000105D55400AA082A8215",
INIT_25 => X"145F7840000000000000000000000000000000000000000000002AB45555568A",
INIT_26 => X"50AAF7F1FDE38FF8A2DA101C2AAFA00EB8E0516DE3F5C000014041256DEBA487",
INIT_27 => X"2FB551C0E0516D417FEDA921C000017DEBF5FDE92080E000BAF7DB4016DE3DF4",
INIT_28 => X"0070BAAAAAADBD70820801EF085F7AF6D55556AA381C75EABEFBED1575C7E380",
INIT_29 => X"DF7AE82F7AA870AA0071F8FFFBE842DA101C0E2DB55410A3FFC7F7A087000FF8",
INIT_2A => X"7DF7DFD7A2A480000BE8A17482F78A28A92E3841556DA2FBD7545F7AAAFABAFF",
INIT_2B => X"41554508208208017DF7F5FDE9208556FBC7A2DB400824120ADA38E3F1EFA28F",
INIT_2C => X"000002DB455D5B68A28A2FFC20AAEB842DAAAE38A02082E3FBC217D1C0E05000",
INIT_2D => X"005504001FFAA8015545F7800000000000000000000000000000000000000000",
INIT_2E => X"0BAFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE10552EBDE00AAAE975FFAAD1420",
INIT_2F => X"8BEFF7D157555AA803DF45552E975EF007FFFE005504001FFAAD17DE00082E82",
INIT_30 => X"BFF55FF8017410FF84154BAAAAABFF450000021FF007BE8BFF5D516AABA5D556",
INIT_31 => X"BD5555F7AEBFEBAFFFBEAA00F7AE974BA085568BEFF7803FE10552EBDF45002E",
INIT_32 => X"003DEAAA2D57FEAAF7FBFDF45AA8002000FFAE95400F7AEA8A10A284175FFAAF",
INIT_33 => X"2FFC21EF552A954100851554000004021FFFFD17DE1008517DF55A2FBC201008",
INIT_34 => X"00000000000000000000003DF55557FEAAAAA2FFC00AAAA803FEAAA2AA82000A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00020201926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"00104884880A4400403000004800027102A0E88110D83210642EA809C0203040",
INIT_05 => X"04092A08138041184109C001380000201A008128044E00754010C9C192D82400",
INIT_06 => X"201800012372A1D72A180000204024024954A3670819290951001009092C0222",
INIT_07 => X"4000220B40020C80052C0A12292A040005715540015E006810001C4B01032C7E",
INIT_08 => X"9032881000140140024200808839005C002010800000155F8122851320016400",
INIT_09 => X"2C80080200801280825A988008000040008208401005B3071859006442004054",
INIT_0A => X"200810940400720005C0030192072310200028B6022346080802E001A5600801",
INIT_0B => X"206822F20CA8826AC2A14250A128509528954404144C200425010040000001B0",
INIT_0C => X"A41AA5B7344C10B383081BA4B7341C10B3831034081200000000000430003000",
INIT_0D => X"381BA4B7344C10B383081AA5B7341C10B383110218CB0E54C2EA404A4F03D404",
INIT_0E => X"A008E730A01AB113A5524E6ACA678001CE3E20A5B284ED1132909C72885A2B2C",
INIT_0F => X"6430202021252991C22C99731014AC3CC0C0B8182597A801610218CB0C3548B3",
INIT_10 => X"5194332B018A444AEA2701288A15A151EC5952E44128CA194517354C180A3C06",
INIT_11 => X"D50048A411C158BB0A7910142C771804C8A0ADA2E6A983014780CA28B2A5C882",
INIT_12 => X"F8BE8E3E1E0109472C3EB50158BB02D09852745F80112C428562EE0353635232",
INIT_13 => X"02414032646000826080C20001104240480068001C9B9150A0000297046E4023",
INIT_14 => X"4510008241C80290882400908000A000A1000809A93485D61000000000000080",
INIT_15 => X"00000000040000000000000020000000000000008010102A82014100101118BA",
INIT_16 => X"A10441010090480C096420184321040002844840000000004000000000400000",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094246A10",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"0000000000005094250942509425094250942509425094250942509425094250",
INIT_1A => X"BFBFBFBF7DDF3BAAAAAABEFDDFE7EFBEFFE7CFC3F7EFFF7DF7E24502A8000000",
INIT_1B => X"F5FAFD7EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAFFD",
INIT_1C => X"BF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EB",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800FFDFAFD7E",
INIT_1E => X"80155F7842AB55552E821FFFFD5555EF552ABDFEF007FE8A00AAFBC000000000",
INIT_1F => X"BD55EFAAD1554BA00556AA00AAD16AA10FF8002155F7FFC2000080417555FFAA",
INIT_20 => X"55420AAF7D542155F7D1400AAF7FFFDE00F7842AA00002A821EF5D7BC21FFFFF",
INIT_21 => X"80000155F7FFFDEAA00002AB45082A821EF5D557FF45A2AABFEBA082A975555D",
INIT_22 => X"A2FFE8BEF5D517FF455D554214500043DEBAAAFFEAB55080000145557FE8AAA0",
INIT_23 => X"0552EBFEAAAAD1401FF08557DF4555516AA00007BEABEFAAD1555FFF7842AABA",
INIT_24 => X"FFFFAE82000FF80020AAA2AAAABFF002E80000AAAABDF555D2E955EFA28428A1",
INIT_25 => X"A28AAF5C0000000000000000000000000000000000000000000028B4555043DF",
INIT_26 => X"000014041256DEBA487145F78428B6D4120851FFEBD5525C74124B8FC71C71EF",
INIT_27 => X"871C74975C01FFEBF5D25EFA2D555482085F6FA28AAD16FA00EB8E0516DE3F5C",
INIT_28 => X"0BFE921C2E9557D415B400BAF7DB4016DE3DF450AAF7F1FDE38FF8A2DA101C2A",
INIT_29 => X"0E0516D417FEDA921C000017DEBF5FDE92080E2AB7D1C24851FF495F7FF55A2A",
INIT_2A => X"ED1575C7E38028A82B6F1E8BFF495F78F7D49554214508003FEAABEFFEFB551C",
INIT_2B => X"5D20905C7AA842DA00492EBFEAABED1401EF085F7AF6D55556AA381C75EABEFB",
INIT_2C => X"000002DB55410A3FFC7F7A087000FF80070BAAAAAADBD7082087000AAA4BFF7D",
INIT_2D => X"4508042AB455D517DEBAA2D54000000000000000000000000000000000000000",
INIT_2E => X"E00AAAE975FFAAD1420005504001FFAA8015545F78028BFF0004175EFA2D5421",
INIT_2F => X"DEAAF7AABDE10552E975450051401EFA2D5421EFAAD557410007BFDEAAA2D57D",
INIT_30 => X"175FF087BFFF45AA843FE005D2A955FF087BC20BAFFFBC01EFA2FFD74AAF7D57",
INIT_31 => X"03FEBAFFFBFDF45552E975EF007FFFE005504001FFAAD17DE00082EA8BFF5504",
INIT_32 => X"516AABA5D5568BEFF7D157555AA8028A00FFD16ABFF087BEABEF005542155000",
INIT_33 => X"00017410AA803DFEF550402155A2843FE00082ABFEAAFFD5421FF007BE8BFF5D",
INIT_34 => X"00000000000000000000003DF45002EBFF55FF8017410FF84154BAAAAABFF450",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000033FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"0002074F200904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000480488024000403000000000001002A0E881108032100002000800203040",
INIT_05 => X"04092A081000411841080001000000201000012800400010001081C000402000",
INIT_06 => X"80500001221021C1021800002000240249048361001128081100100909000222",
INIT_07 => X"4000220050020480152D0A142D0A8400043B45400040006810000C5901033D78",
INIT_08 => X"0010880000100140024280808829029C002000000000053FA142051324902030",
INIT_09 => X"2000000000000200820888800800004000800840100020011858006442004040",
INIT_0A => X"200800840400400005C0010190070310200008B202236D080802400001600801",
INIT_0B => X"000000100C088020028102408120409120940404104C20002101004000000110",
INIT_0C => X"5210040000B0E0A0000210040000E0E0A0000190081200000000000000003000",
INIT_0D => X"0210008000B0E0A0000210008000E0E0A0000B02740421A0E5D1A02400205080",
INIT_0E => X"40110080A4006110510C14D18178E01200860008920106460D4501CB00011130",
INIT_0F => X"411420220080220C0093C38923240ABBC00905C33C6000400F02740412C0715C",
INIT_10 => X"8000120800658992F3C700C3018120000041DB011CC000090012565306500002",
INIT_11 => X"E240240A8340000200067EAA8CB65809240C09024A4AE0CA0000480083968239",
INIT_12 => X"7DB0D0200900422ACA4B28000002002B46867DBC002A830280000800F7B7A0B1",
INIT_13 => X"020040126060008020000200000042004005800004801150A00341244000845C",
INIT_14 => X"4500008240800000802000908000800001000009A92481041000000000000080",
INIT_15 => X"000040000000000000040000000000000000000080101000000141001001088A",
INIT_16 => X"810440000090480C096420084101040000044040000000004000040000000000",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090246810",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"0000000000004090240902409024090240902409024090240902409024090240",
INIT_1A => X"EFBBBBAABCDABF9E79E7BEF9CB91FE1EF7D3AEB9F3E6FF7DF650400280000000",
INIT_1B => X"FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7FC",
INIT_1C => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8FF000FE7F3F",
INIT_1E => X"E8A00AAFBE8BEFA2D568ABA00003DF555555574AAAAAEAAB45082E8000000000",
INIT_1F => X"02AABA555155400557BC2010557BEAB55552E821FFFFD5555EF552ABDFEF007F",
INIT_20 => X"002AA10FF8002155F7FFC2000080417555FFAA80155F78428AAA007FE8A10080",
INIT_21 => X"AD1554BA00556AA00AAD140145AA8028ABA002EBFFFF082EBDEBAA2D1420105D",
INIT_22 => X"A2AEA8A10080428A10FFAEBFFEF5D0428B45A2FFC21EF5D7BC21FFFFFBD55EFA",
INIT_23 => X"5F7FBC0010FFAA820AAF7D542155F7D1400AAF7FFFDE00F7842AA00002A80155",
INIT_24 => X"EF5D557FF45A2AABFEBA082A975555D55400BA005568A000000175FFF7D15554",
INIT_25 => X"B6D00248000000000000000000000000000000000000000000002AB45082A821",
INIT_26 => X"25C74124B8FC71C71EFA28AAF5E8BFFB6D56DA82000E38F6D4155504AAA2AEAA",
INIT_27 => X"28ABA147FEDA10080E2AAAA555552400417FC20005D75E8B6D4120851FFEBD55",
INIT_28 => X"4BAEAAB6DB4202849042FA00EB8E0516DE3F5C000014041256DEBA487145F784",
INIT_29 => X"75C01FFEBF5D25EFA2D555482085F6FA28AAD147155BE8028A82002EB8FC7002",
INIT_2A => X"F8A2DA101C2A80145B6AEA8A10080E2DA00F7A0BDFD7550428B55A2F1C71C749",
INIT_2B => X"0004175FFE3D15757DE3F5C0038FFAA800BAF7DB4016DE3DF450AAF7F1FDE38F",
INIT_2C => X"000002AB7D1C24851FF495F7FF55A2A0BFE921C2E9557D415B400AA00556DA00",
INIT_2D => X"EF0051400AAA2AAAABFF08000000000000000000000000000000000000000000",
INIT_2E => X"BFF0004175EFA2D54214508042AB455D517DEBAA2D568BEFFFD57FE10002AAAB",
INIT_2F => X"01FFAA8015545F78028AAA557FFFE00082EAAAAA5D5142000007BC20105D5568",
INIT_30 => X"28A00082EAAB45000028ABAFFFBC20AA08043DE00AAAE975FFAAD14200055040",
INIT_31 => X"02AB55AAD1575450051401EFA2D5421EFAAD557410007BFDEAAA2D557555FF80",
INIT_32 => X"FFD74AAF7D57DEAAF7AABDE10552E82155FFAAA8A10002ABFE00F7803FF555D0",
INIT_33 => X"87BC20AA00517DE000804175EFAAD1555EFA2D1420BAFFAE820BAFFFBC01EFA2",
INIT_34 => X"000000000000000000000028BFF5504175FF087BFFF45AA843FE005D2A955FF0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000100000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"000440009282000001100000000000100220C8811080321000000228002A3000",
INIT_05 => X"04092A0010004300418800510000A6201000012A64400000145080C000422000",
INIT_06 => X"00100001220001C00018821020402402080003772019200001001009090002AA",
INIT_07 => X"4000220000021840010C8912250A0400042044400040006810000C4901032B18",
INIT_08 => X"0022810000058140024280A0A8190004002030C00000016F8122041320000000",
INIT_09 => X"20000000000002C0820888008800000000800840100020011850004402004040",
INIT_0A => X"00080094000062000180010180060210200008B2022304080800400003E00801",
INIT_0B => X"0000000008008020020000000000000100800000000000002500004000000130",
INIT_0C => X"0010108000000000000010108000000000000230001200000000000420003000",
INIT_0D => X"0010140000000000000010140000000000000100000040000000000000000000",
INIT_0E => X"0000000000000100008040000000000000000000020000090000000000000000",
INIT_0F => X"0030002000406000000000068409014000000000000000000100000040000000",
INIT_10 => X"0000000800000201000800000000000000400048000000000010000440000000",
INIT_11 => X"00A0000000000002000000441108800000000002008008000000000080201000",
INIT_12 => X"0242038B82800000000000000002000001000000000000000000080000001844",
INIT_13 => X"000000100000000005C04A000000400000000000000001062000000400000000",
INIT_14 => X"4500008200800000800000100000800001000001A12480001000000000000080",
INIT_15 => X"000000000000000000040000200002000000000080101000004140001001088A",
INIT_16 => X"0004400000904808094020080000000000044040000000004000040000400004",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000046000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000400280000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000000000",
INIT_1E => X"AAB45082EBFE000004020AA552E80000F7FBC214555003DE10A2FBC000000000",
INIT_1F => X"BE8A10F7802AA0055003FE10007BE8BEFA2D568ABA00003DF555555574AAAAAE",
INIT_20 => X"AEAAB55552E821FFFFD5555EF552ABDFEF007FE8A00AAFBFDEBA555568BEFA2F",
INIT_21 => X"55155400557BC2010557BFFFEFA2FFC20005D2A955EFF78428BEFAAD17DF55AA",
INIT_22 => X"5D2AA8B45AAD57FF55A2FBC21FFA28415400FF8028AAA007FE8A1008002AABA5",
INIT_23 => X"A002E9740055516AA10FF8002155F7FFC2000080417555FFAA80155F7843DF45",
INIT_24 => X"BA002EBFFFF082EBDEBAA2D1420105D003FFFF08514200055002AA00AA802AAB",
INIT_25 => X"E28B6FFC0000000000000000000000000000000000000000000000145AA8028A",
INIT_26 => X"8F6D4155504AAA2AEAAB6D0024B8E381C0A00092412A87010E3F5C0145410E3D",
INIT_27 => X"F8EAA495F68BFFA2F1EFA38E38428A005D0038E28147FE8BFFB6D56DA82000E3",
INIT_28 => X"428BEFB6DB7DF45AAAEA8B6D4120851FFEBD5525C74124B8FC71C71EFA28AAF5",
INIT_29 => X"7FEDA10080E2AAAA555552400417FC20005D75F8FFFBEF5C0000492A955FFF78",
INIT_2A => X"BA487145F7843FF7D4120A8B6DAAD17FF55B6F5C21EFAA8E10400E38E28ABA14",
INIT_2B => X"41002FA38A2842AA82142095428415F6FA00EB8E0516DE3F5C000014041256DE",
INIT_2C => X"0000007155BE8028A82002EB8FC70024BAEAAB6DB4202849043FFC7005F45010",
INIT_2D => X"00A2D542155002ABDEBAF7FBC000000000000000000000000000000000000000",
INIT_2E => X"BEFFFD57FE10002AAABEF0051400AAA2AAAABFF08002AAAA5D2A82000082E954",
INIT_2F => X"AB455D517DEBAA2D56AABA087BEABEFAAD57DEAAA2802AA105D002AABA5D7BE8",
INIT_30 => X"42010082A955EFFF8428BFFFFFBFDF55A2AEA8BFF0004175EFA2D54214508042",
INIT_31 => X"A82000AAAAA8AAA557FFFE00082EAAAAA5D5142000007BC20105D556ABFFF7D1",
INIT_32 => X"D1420005504001FFAA8015545F7803FFEF08002ABEFA2D57DF45F7D1401FFA2A",
INIT_33 => X"8043FF55087BD740000043DEAAA2842AA005D00154AA007BFDE00AAAE975FFAA",
INIT_34 => X"000000000000000000000017555FF8028A00082EAAB45000028ABAFFFBC20AA0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000300000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"0202115002BB10080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"2FE962000017102918900948514522CE09200C0D590569398ADBF8CC1E50E480",
INIT_05 => X"5E6023002834854AE41C1E8782F508F2A15B71D412E0AFD9C2990DA56FF0B55A",
INIT_06 => X"B9B9E55402000340003200220A86012D0000000480D0400001555960540180A0",
INIT_07 => X"40D890101DBD400901442800817C2901F400868554DE240000A80090CE82A803",
INIT_08 => X"0122004000005665510320C9C90510025A8A00000A0A048F550A440E0001380C",
INIT_09 => X"2060410280081116C8204D016CB2CB290008008279580411289000000118A905",
INIT_0A => X"00008176802203180025699200140001A15000017F0051D0F837324E002A8A56",
INIT_0B => X"4485D000000124002400000000000001004010A8812831605DA0000A054052E4",
INIT_0C => X"B5320018CAC99BA0A3B9320018CAAAADA0C343F1AC1B01040A00202489551455",
INIT_0D => X"59320018CAC99BA0ACB9320018CAAAADA0CC421CA003B694B68018FAAA708E2C",
INIT_0E => X"B2449A3FF2FA04E5E09B128834ADB1443A1891E4A928C29020E6A8524CE7A3EE",
INIT_0F => X"2375B801324301AB0067622E5E5404B2A5A40B1E6644AF0F021EA003AC24352A",
INIT_10 => X"0A8C241815FEB6A9158863F638FB60ED838E890B703C6260D8E3A21275714C90",
INIT_11 => X"15F11133D171727A2550EE2F1BA0064F70DBDB1C74424E91E1C194C71D1216F5",
INIT_12 => X"432A2B2D001F803471A9A960E57245FDF9D364DBD9435A6D45C9E81BED555E4C",
INIT_13 => X"C00006B0800000038814B72AB01508150013F162119014204373517700ACCC59",
INIT_14 => X"300208092B940192D1000000000000A8A5AA80018120E00066000000000012CA",
INIT_15 => X"1000110001100011000108000880008000520228080108039501200848002912",
INIT_16 => X"081500008A422150884081AC9000010003561180063DB4F61100011000110001",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000012000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"BCBF0F2C688A8D3CF3CF0A7A898D21B4C9838D3030EF5168A360400000000000",
INIT_1B => X"E9F47A7D345345345345345345345345345345345345345145145145145147A5",
INIT_1C => X"3E9F4FA3D1E8F47A3D1E8F47A3D1E9F4FA7D3E9F4FA7D3E9F4FA7D1E9F47A7D1",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800001F4FA7D",
INIT_1E => X"3DE10A2FBC21FFFFFBFDF45A2D56AB45FFFFD54BAFF80001FF002A8000000000",
INIT_1F => X"FFFE005D7BC0010002E954AA087FFFE000004020AA552E80000F7FBC21455500",
INIT_20 => X"FFE8BEFA2D568ABA00003DF555555574AAAAAEAAB45082E974BA5D7BFDF55A2F",
INIT_21 => X"7802AA0055003FE10007BC0000082A97400550017410FFD1555550000020BAAA",
INIT_22 => X"AAFBD74105504021FF5D2EAAABAFFFBD55FF002ABDEBA555568BEFA2FBE8A10F",
INIT_23 => X"0007FC00AA087FEAB55552E821FFFFD5555EF552ABDFEF007FE8A00AAFBD55EF",
INIT_24 => X"005D2A955EFF78428BEFAAD17DF55AAAE820AA5D517DF45AAFFFFEAAFFAABFE1",
INIT_25 => X"1FF08248000000000000000000000000000000000000000000003FFEFA2FFC20",
INIT_26 => X"7010E3F5C0145410E3DE28B6FFC21C7E3F1F8F55AADB6FB6DFFFBD54AAE38E02",
INIT_27 => X"92482497BFDF45AAFFF8E385D7BC5000002E904BA1C7FF8E381C0A00092412A8",
INIT_28 => X"B555450804070BABEF5E8BFFB6D56DA82000E38F6D4155504AAA2AEAAB6D0024",
INIT_29 => X"5F68BFFA2F1EFA38E38428A005D0038E28147FC2010142E90428490015400FFD",
INIT_2A => X"C71EFA28AAF5D25D7B6F1D54384904021FF5D2AADAAAFFF1D55FF002EB8EAA49",
INIT_2B => X"A2F1FDEAAEBAABDE001471C20921475E8B6D4120851FFEBD5525C74124B8FC71",
INIT_2C => X"0000038FFFBEF5C0000492A955FFF78428BEFB6DB7DF45AAAE820925D5B7DF45",
INIT_2D => X"EFF7FFD54AAAAAA801EF00000000000000000000000000000000000000000000",
INIT_2E => X"AAA5D2A82000082E95400A2D542155002ABDEBAF7FBC2145AAD568B45AAFBFFF",
INIT_2F => X"00AAA2AAAABFF080000000087BFDF55A2FFE8AAA557FD7410082A800AA557BEA",
INIT_30 => X"800BA080417400F7FBD75450800174AAFFD168BEFFFD57FE10002AAABEF00514",
INIT_31 => X"1575EF082EAAABA087BEABEFAAD57DEAAA2802AA105D002AABA5D7BC20005D2E",
INIT_32 => X"D54214508042AB455D517DEBAA2D540155F7D1554AA0800001EF5D2ABDEBAF7D",
INIT_33 => X"2AE82010557FFDF55A2D57FEAAAAAEBFE10555140000555568BFF0004175EFA2",
INIT_34 => X"00000000000000000000002ABFFF7D142010082A955EFFF8428BFFFFFBFDF55A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000100000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"5295B6957FCBE0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"6DE90201BF90102103AF158E805428249851BFB2C106592088DBF8400A5055C2",
INIT_05 => X"3824BD7F80148D9E07100A8201ED01C1A19B68F40A807ED9C18114956FF081DB",
INIT_06 => X"6A8F033DD800000000050716BE9F57F8AC000807DFD9B00000CF20E5E1818B1B",
INIT_07 => X"86481240FE05A109228E2C0891D772A6F40045B8CF30E085DD2ED57D4EED08CA",
INIT_08 => X"DF23800005981C0338190549C904182B6113870022000488C08B46268A001508",
INIT_09 => X"823DF78CDB6CA60E0E28EFFE2061872F80C1684A80C8604085F0074D3B72637F",
INIT_0A => X"BD2FAD7FE653C3BA1FF33E0E001E000B3A5DAADAFDDA5DA79350CFB8013E7437",
INIT_0B => X"C5C3D00018006C681700000000000000020012E9E10A31EB5FF9296A67F5B4FF",
INIT_0C => X"542A6FEEB2533EA160782A6FEEB2333EA16031F2BD47BDA2CA5D8164FCCFE833",
INIT_0D => X"F82A6FEEB2533EA160782A6FEEB2333EA160391BEFF2C32FB695F919110D5ECE",
INIT_0E => X"5A86840354D1706FFFA3EF6E24B6D18C0D06638A207CFDE1F7DDAD76D5282400",
INIT_0F => X"4D77FAAB77CE3AF3EE78F58DB737E6E43E59AFE4A59B57679D19EFF2C7573FAD",
INIT_10 => X"72CA52606DFED6CA55334C04C04FF7D7A0ABD6DAAAB96529382B74E4E1FE4ACA",
INIT_11 => X"AA1A184045D5D7A870D2F5A5D7522D1281017F056E9C9C3FC95949C157ADB555",
INIT_12 => X"A58949D5B5C85F97871876F7D7E859FDEB974F486905001FDF5FA0D719F9956E",
INIT_13 => X"70021EE341036BF368128419FB5560158015177F916A039EF41FDB34A91F432E",
INIT_14 => X"1D0A7CC9AE7A08BFF0001D35682AC0CE8FCCC200A59BDD2FFE3F3EC7C7DEF206",
INIT_15 => X"BCF4FBCF4FBCF4FBCF4FBE7A7DE7A7800617112E46F05D02DD814102F800633F",
INIT_16 => X"00179C16DECF67F08BC02F9086000D9E8A3F06ABD73DBCF4FBCF4FBCF4FBCF4F",
INIT_17 => X"000000000000000000000000000000000000000000000000000000000005F080",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"930D0D1B9000303AEBAE88BE013DB9880A5D25C0408006114F981800C0000000",
INIT_1B => X"351A8D069A6BAE9A69A6BAE9A6BAE9A69A6BAE9A6BAE9A69A69A69A69A69A918",
INIT_1C => X"A351A8D46A351A8D46A351A8D46A341A0D068341A0D068341A0D068351A8D068",
INIT_1D => X"00000000000000000000000000000000000003FFFFFFFFFFFFFF8000011A8D46",
INIT_1E => X"001FF002A821FFFFFFFFFFFFFFBFDFEFAAD142010007BEAB55FFAA8000000000",
INIT_1F => X"A975EFA2D140145007BC21FF5D2A821FFFFFBFDF45A2D56AB45FFFFD54BAFF80",
INIT_20 => X"7BFFE000004020AA552E80000F7FBC214555003DE10A2FBEAB45A28000010082",
INIT_21 => X"D7BC0010002E954AA087FD7400082E954AA0800154AA0855575FFAAD57FE005D",
INIT_22 => X"F7D16AB45FFFFEABEF007BD74005555555EFF7AE974BA5D7BFDF55A2FFFFE005",
INIT_23 => X"5555568B45552EA8BEFA2D568ABA00003DF555555574AAAAAEAAB45082EBFFFF",
INIT_24 => X"00550017410FFD1555550000020BAAAFFC0145AA84154BA082E801FFAAFBC015",
INIT_25 => X"B7DEBA480000000000000000000000000000000000000000000000000082A974",
INIT_26 => X"FB6DFFFBD54AAE38E021FF0824851FFFFFFFFFEFF7F1FAFD7A2D5400001C7BED",
INIT_27 => X"EFB45AA8E070281C20925FFBEDB451451C7BC01EF4124821C7E3F1F8F55AADB6",
INIT_28 => X"5505EFBEDB7AE385D7FF8E381C0A00092412A87010E3F5C0145410E3DE28B6FF",
INIT_29 => X"7BFDF45AAFFF8E385D7BC5000002E904BA1C7FD54280024924AA1404174AA005",
INIT_2A => X"2AEAAB6D0024BFFD7FFDB6AB7DFFF5EDBC71C7BD54005D5B575EFEBAE9248249",
INIT_2B => X"1C20801FFB6F5C0145555B68B7D4124A8BFFB6D56DA82000E38F6D4155504AAA",
INIT_2C => X"0000002010142E90428490015400FFDB555450804070BABEF5C516DAA8A12492",
INIT_2D => X"45AAD5400005D7BFFFEFAA800000000000000000000000000000000000000000",
INIT_2E => X"145AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF0000155FFF7FBFDFEFFFD568B",
INIT_2F => X"2155002ABDEBAF7FBFDF55A2AA974AA5D04001EFFFFFD5545557BC21FF080002",
INIT_30 => X"000AA5500174AA0855421FFFFFBEAAAA5D7BEAAAA5D2A82000082E95400A2D54",
INIT_31 => X"BD75FFAAAA80000087BFDF55A2FFE8AAA557FD7410082A800AA557BD74BA0004",
INIT_32 => X"2AAABEF0051400AAA2AAAABFF08003FF55F7FFEABFFF7D57FF455D7FD54105D7",
INIT_33 => X"FD1555FFA2AA800105504001EFFFD140145557BE8BEF000028BEFFFD57FE1000",
INIT_34 => X"0000000000000000000000020005D2E800BA080417400F7FBD75450800174AAF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000033FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"080BA868803F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"42016B0C401F58495C900A4859552A611D9A640F5903B2388004004C08A06008",
INIT_05 => X"16226B107811422A641C08038040007060E0032801E0202000991B708280B501",
INIT_06 => X"B3B8E0FC86142B4142B0000000011114D305824024090A1A143F182000000000",
INIT_07 => X"802102401015610A02C4005000EA019D002482043FCF1C8090C02800C0120886",
INIT_08 => X"20D40A5004003260F9810541494D403D9B98810A0002C601000054B94A006880",
INIT_09 => X"6070000504102805C820C8016C30C250080C0182183804012A0A102200110180",
INIT_0A => X"E000108010230445A800FD865421432121804021C20452880C2D100000022E0C",
INIT_0B => X"C2060014250B9080008306C18360C1B0609C05013065CC042004040808084001",
INIT_0C => X"8582081483ACC15F9C3982081483CCC15F9CBA45505640000A402019003F140F",
INIT_0D => X"F982081483ACC15F9F3982081483CCC15F9FB1962FCB69E08AAAEAEBCDDF7C72",
INIT_0E => X"E3F8E7F5E3AC3620805298B15A3FEBF1CFFF7670ACC3811A28AB57523CDFEBFB",
INIT_0F => X"DC4041D4CF03138DD865103EFEEAC9002BF05800D875E63CC9962FCB52CAA02F",
INIT_10 => X"8DB7BFE25208E8F46A228BF8A757F1B72A8A800B7546DB9F1CA320037F01BD67",
INIT_11 => X"9509EAAE7FD3B749471C48F8A45981CCFAFDBF9464006FD037AEFAE5150016EA",
INIT_12 => X"8802A3AF8E8FB0440CE78773B709641256EC844B8AF92FD7CEDC24A9E181A8A2",
INIT_13 => X"C284601C2864000080113307E4800297D086E00036D2440E0880AAD62BEFF577",
INIT_14 => X"A88DCC2211E44174112840880000060D7030C30B885200D274004008080003C1",
INIT_15 => X"0308003080030800308001840018400400602A01880980037109700C04C44C92",
INIT_16 => X"8340000020301805002D008CD943626111C0D95C20C2030A0030800308003080",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B0680834",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"00000000000041B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1",
INIT_1A => X"60B22A145DF60B8208209679D701DC2E784601F95163897DF160000000000000",
INIT_1B => X"944A2512AAA8A28A28A2AAAAAA8A28A28A2AAAAAA8A28A28A28A28A28A28A244",
INIT_1C => X"8944A25128944A25128944A25128944A25128944A25128944A25128954AA552A",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8000004A2512",
INIT_1E => X"EAB55FFAA821FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E820BA55000000000000",
INIT_1F => X"16AB55A2D542000A2D5400BA0800021FFFFFFFFFFFFFFBFDFEFAAD142010007B",
INIT_20 => X"80021FFFFFBFDF45A2D56AB45FFFFD54BAFF80001FF002A821FFFFFFFFFEFF7D",
INIT_21 => X"2D140145007BC21FF5D2AAABFFF7D168B45AAD57DFFFFFFFC0010F7842AA10F7",
INIT_22 => X"000002010552E95410AAFBD75FF5D7FEAB5500516AB45A28000010082A975EFA",
INIT_23 => X"5A284155FF5D517FE000004020AA552E80000F7FBC214555003DE10A2FBEAA00",
INIT_24 => X"AA0800154AA0855575FFAAD57FE005D7BD74000804174AA5D00020BA55554214",
INIT_25 => X"0AA490A00000000000000000000000000000000000000000000017400082E954",
INIT_26 => X"AFD7A2D5400001C7BEDB7DEBA4871FFFFFFFFFFFFFFFFDFEFF7FFD74AA552A82",
INIT_27 => X"821FFF7F1F8FC7EBD568B7DB6DF47000AADF400AA080A051FFFFFFFFFEFF7F1F",
INIT_28 => X"1C2000F78A2DA38E38A021C7E3F1F8F55AADB6FB6DFFFBD54AAE38E021FF0824",
INIT_29 => X"8E070281C20925FFBEDB451451C7BC01EF4124ADBC7E3D56AB7DB6DF78FD7EBF",
INIT_2A => X"10E3DE28B6FFE8A101C0E05010412495428AAF1D25EF497FEAB7D145B6FB45AA",
INIT_2B => X"5D0A000BA555F47145BE8A105EF555178E381C0A00092412A87010E3F5C01454",
INIT_2C => X"00000154280024924AA1404174AA0055505EFBEDB7AE385D7FD7438140012482",
INIT_2D => X"EFFFFBD54BA5D2A820AA082A8000000000000000000000000000000000000000",
INIT_2E => X"5FFF7FBFDFEFFFD568B45AAD5400005D7BFFFEFAA80155FFFFFFFFFFFF7FBFDF",
INIT_2F => X"54AAAAAA801EF0000021EFF7D16AB55A2D56ABEFF7FBD5410AAFBC00AA002A95",
INIT_30 => X"68BFFF7FFEAB45AAD140010F7AABFEBAAAAA82145AAD568B45AAFBFFFEFF7FFD",
INIT_31 => X"BE8BFF557BFDF55A2AA974AA5D04001EFFFFFD5545557BC21FF08003FF55AAD1",
INIT_32 => X"2E95400A2D542155002ABDEBAF7FBE8A00552E954100000154AAA2D1421FF007",
INIT_33 => X"D7BD74BA5D0002010552E820AA5D7BD7545F7AA801EF55516AAAA5D2A8200008",
INIT_34 => X"0000000000000000000000174BA0004000AA5500174AA0855421FFFFFBEAAAA5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000100000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000010228001000000000000000000024001620280000000000354200004008",
INIT_04 => X"00016200001310090090004840004152C7208802590000388000004C08006000",
INIT_05 => X"1621008008100002641C0803804000702000000000E02000009900000000B100",
INIT_06 => X"0210200C00000000000000000000000080000000000000000003182000000000",
INIT_07 => X"C00D267001B880080700285020020AC98820022802400480405008901100A001",
INIT_08 => X"000000000000106009872048400C4000010D000008000204150A00815A010084",
INIT_09 => X"0000000000000004C80000002C30C200000000021808005800000000000E0E00",
INIT_0A => X"0000000000000000080025860000000080A00020602040800000000000022A04",
INIT_0B => X"C002000000000000000000000000000000000000000000000000000084000760",
INIT_0C => X"385598035D0008A003B05598035D0008A0034078104B41A41000000000031400",
INIT_0D => X"505598035D0008A000B05598035D0008A0004263C0343EDD414004042228DC0D",
INIT_0E => X"0401180DE053A98F6ECC739D8140040231068187C39F5A4F985C008902041124",
INIT_0F => X"227848D4303807FC8CC5508AEAED1BFBD406451B02000E033263C0343CB74050",
INIT_10 => X"00000018A700FCF980CC300318A2420851546B2400000040D8549B5800000010",
INIT_11 => X"40E40511802208D6B30C48F8A8A452210402120A936B0000000004C2A8D64800",
INIT_12 => X"0006362A2B6424287B08286208D6B1427ED430B41402D025082359700181C211",
INIT_13 => X"40000000000000000010030060009C000018440021011821B35254E99AF9E941",
INIT_14 => X"002000044000000000000000000002F0001F00002024B20002000000000002C0",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000040",
INIT_16 => X"00000000000000000000008C8000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"441189B9045D82A69A69803F47E18E0218CC0140400200441920000000000000",
INIT_1B => X"4C261309861861861A69861861861861A69861861861861861861861861861A1",
INIT_1C => X"84C26130984C26130984C26130984C26130984C26130984C261349A4C2613098",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000261309",
INIT_1E => X"820BA55003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A800105D2E8000000000",
INIT_1F => X"FFDFEFF7FFD54BA5D2EA8BFFFF84021FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E",
INIT_20 => X"AE821FFFFFFFFFFFFFFBFDFEFAAD142010007BEAB55FFAABDFFFFFFFFFFFFFFF",
INIT_21 => X"2D542000A2D5400BA08003DFFFFFFFFFFFFF7FBE8B55A2D540010007BEAABAA2",
INIT_22 => X"FFFFFDFEFA2D56AB45AAFBD74AAFFD5420100804021FFFFFFFFFEFF7D16AB55A",
INIT_23 => X"AFF802ABFFFFAE821FFFFFBFDF45A2D56AB45FFFFD54BAFF80001FF002ABDFFF",
INIT_24 => X"45AAD57DFFFFFFFC0010F7842AA10F780155FFF7FBE8B45AAD568BFFF7FBD74B",
INIT_25 => X"000412A8000000000000000000000000000000000000000000002ABFFF7D168B",
INIT_26 => X"DFEFF7FFD74AA552A820AA490A38FFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2A80",
INIT_27 => X"BAFFFFFFFFFFFFF7FBFDFD7EBF1D24AA5D2AADBD7E384071FFFFFFFFFFFFFFFF",
INIT_28 => X"140000007FEFA92A2AA851FFFFFFFFFEFF7F1FAFD7A2D5400001C7BEDB7DEBA4",
INIT_29 => X"F1F8FC7EBD568B7DB6DF47000AADF400AA080A3FFFFFFFBFDFC7E3F5EAB45AAD",
INIT_2A => X"38E021FF0824BDFEFE3F1F8FD7AAD16DB7DBEFBD74AAE3DF400000004021FFF7",
INIT_2B => X"B6DB6FBD7E3F5D04AAFF8A2DBD7E3A0821C7E3F1F8F55AADB6FB6DFFFBD54AAE",
INIT_2C => X"000002DBC7E3D56AB7DB6DF78FD7EBF1C2000F78A2DA38E38A125C7E3F1EAB55",
INIT_2D => X"FFF7FBD54BA552A80010002A8000000000000000000000000000000000000000",
INIT_2E => X"5FFFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA082AA8BFFFFFFFFFFFFFFFFFF",
INIT_2F => X"00005D7BFFFEFAA8028BFFFFFFFDFEFF7FFFFF55A2D5400AA552ABDF55A28015",
INIT_30 => X"FDF55AAD16AB55AAD140010007BFFE10AAAA955FFF7FBFDFEFFFD568B45AAD54",
INIT_31 => X"BC20100800021EFF7D16AB55A2D56ABEFF7FBD5410AAFBC00AA002ABDFEFF7FB",
INIT_32 => X"FBFFFEFF7FFD54AAAAAA801EF00003FFEFA2D56AB45A2D57DFFFFFFFD54AAA2F",
INIT_33 => X"AAA82155AAD568B55FFFFFDF55A2D1400AAF7AABFF45AA8002145AAD568B45AA",
INIT_34 => X"00000000000000000000003FF55AAD168BFFF7FFEAB45AAD140010F7AABFEBAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000200000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"0001E6000053300B00D0005800000000000000407B0004BB830004DC3D01E000",
INIT_05 => X"FEE0000008720043EC3C3D0F87FA19F7E0201C409BE1F10623BB000A100CF300",
INIT_06 => X"06102FFC8E0007C00078008000171175A200096404D9404003FFDBE4744200AA",
INIT_07 => X"482491301000010001DC00000000000000004203FE4005800000008030002000",
INIT_08 => X"20E2008000027FEFF946058180010429000001080AAA010F8000000000000000",
INIT_09 => X"400000120000913FD80000003DF7DE0080010047FBF8000000000800C5408000",
INIT_0A => X"0080000010000400080FFDBE000000400000010000010050600220461003EAFE",
INIT_0B => X"C00600000000801020000000000000010240001721214E000004000000080000",
INIT_0C => X"08020000200000000F30020000200000000F3008001E00000000001803FF14FF",
INIT_0D => X"F0020000200000000F30020000200000000F3040200000020000000026A70C00",
INIT_0E => X"000019B140000800800000020000000030B86000400080000200000000004A58",
INIT_0F => X"AC08000000508001030A0A4001000000000002183E61E6000040200001000000",
INIT_10 => X"0000A56000090100000000001F86C00010080000000000525801000000000014",
INIT_11 => X"0000001716800000803102020000000002BC360020000000000292C010000000",
INIT_12 => X"DF70C08040100000706707600000801000000000000057450000100106060000",
INIT_13 => X"C011001C81080001101F977FE00800000000000040040040002000080506049C",
INIT_14 => X"0000000000000000020020029000000000000000020000000000000000000ADF",
INIT_15 => X"0000000000000000000000000000000000000000000002000200000000000000",
INIT_16 => X"0801810100000000000093ED8000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000401008080",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"930424038000343CF3CF349600704000201120A983400E0104D2040020000000",
INIT_1B => X"190C86432CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB0C30C30C30C30C818",
INIT_1C => X"2190C86432190C86432190C86432190C86432190C86432190C86432190C86432",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8000010C8643",
INIT_1E => X"800105D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8201008040000000000",
INIT_1F => X"FFFFFFFFFBD54BA552A8001000003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A",
INIT_20 => X"2E821FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E820BA5500001FFFFFFFFFFFFFF",
INIT_21 => X"7FFD54BA5D2EA8BFFFF843FFFFFFFFFFFFFFFFFFFFEFF7FFD74BA552E801FF00",
INIT_22 => X"FFFFFFFFFFFFBFDFEFFFD542000082EAAB55AAAABDFFFFFFFFFFFFFFFFFDFEFF",
INIT_23 => X"0087BE8B55F784021FFFFFFFFFFFFFFBFDFEFAAD142010007BEAB55FFAA801FF",
INIT_24 => X"FFF7FBE8B55A2D540010007BEAABAA2AE975FFFFFFFFFFFF7FBFDF55AAD14000",
INIT_25 => X"00014000000000000000000000000000000000000000000000003DFFFFFFFFFF",
INIT_26 => X"FFFFFFFBD54AA5D2A80000412ABFFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A82",
INIT_27 => X"021FFFFFFFFFFFFFFFFFFEFF7FBD74BA5D2A800281C0038FFFFFFFFFFFFFFFFF",
INIT_28 => X"FD54BA5D2A801C7142E871FFFFFFFFFFFFFFFFDFEFF7FFD74AA552A820AA490A",
INIT_29 => X"FFFFFFFF7FBFDFD7EBF1D24AA5D2AADBD7E38438FFFFFFFFFFFFFFFBFDFEFFFF",
INIT_2A => X"C7BEDB7DEBA4871FFFFFFFFFEFF7FBF8FD7E3D140010142AAFB7DBEAEBAFFFFF",
INIT_2B => X"E3F1FAF45A2D142010087FEDB55F78A051FFFFFFFFFEFF7F1FAFD7A2D5400001",
INIT_2C => X"000003FFFFFFFBFDFC7E3F5EAB45AAD140000007FEFA92A2AA925FFFFFFFDFEF",
INIT_2D => X"FFFFFFD74AA552A820005D040000000000000000000000000000000000000000",
INIT_2E => X"BFFFFFFFFFFFFFFFFFFFFF7FBD54BA552A80010002ABFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"54BA5D2A820AA082A821FFFFFFFFFFFFFFBFDFEFF7FFD74AA5D2A800BA550428",
INIT_30 => X"FFFEFF7FBFFFFFF7FBD74BA552A80145552E955FFFFFFFFFFFF7FBFDFEFFFFBD",
INIT_31 => X"ABFFFFFFAEA8BFFFFFFFDFEFF7FFFFF55A2D5400AA552ABDF55A2802ABFFFFFF",
INIT_32 => X"D568B45AAD5400005D7BFFFEFAA80175FFFFFBFDFEFF7FFEAB45AAD1420105D2",
INIT_33 => X"AAA821EFF7FBFDFFFAAD168B55A2D542010007BFDF55F7AE955FFF7FBFDFEFFF",
INIT_34 => X"00000000000000000000003DFEFF7FBFDF55AAD16AB55AAD140010007BFFE10A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"1094EC681244819000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"0001E6000053300F01D4587800446194F49020107F0012BBC00202DC3823EA82",
INIT_05 => X"FFF201B228704123FC3C381F87C03DFFF012412A9FE1E01013BF09404050F300",
INIT_06 => X"96F43FFF002004020044041084CB01AD000003761702401000FFDFE050000080",
INIT_07 => X"043C802A821D41412001A0040950AB60014114C3FE4187A009A663A680100B30",
INIT_08 => X"2C01004000047EFFF811A46968004060629A0002208A00000068113205A12034",
INIT_09 => X"0A812D8D5B742D3FF84056383FF7DE0880042107BFF9C45B85101C49A37F4000",
INIT_0A => X"0822189000480406310FFDFE00040009814C089202225412115414601DE3EBFE",
INIT_0B => X"C0281280080180B2948004400220011100841200D001000624000100C002804A",
INIT_0C => X"60694101816002D41A4068C101815004D8158809C86065941840B1014FFF56FF",
INIT_0D => X"0068C101816002D41A40694101815004D815810D42E04A08A80098C024500253",
INIT_0E => X"12682960828F05C96A001B029010134160C8125B0B271802242880A04482418A",
INIT_0F => X"100920C54E8EA256ECF078BA081C10080E05C0B06AA8B12CFD0D42E0441A3000",
INIT_10 => X"4F30A8801406D00290006280320100010362A8A20826A88660D86B202049F115",
INIT_11 => X"2011819E290048A2118EC8140C08064802C0081B0D64040936443306C5514410",
INIT_12 => X"C40A0300600C0A80509F418008804581BA0038005A706680012280506A801060",
INIT_13 => X"C000120080002341881F3FFFF80DCC158092C044600466208CC5091011C322A4",
INIT_14 => X"398C6021569249C4B3007127080806FF917FC30010107688862A28C54518DBFF",
INIT_15 => X"228D9228D9228D9228D99146C9146C84006309044081A001B188300E20806520",
INIT_16 => X"8004000000E07008010003EF80022A51904595123203040D9228D9228D9228D9",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010044800",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"0000000000004010040100401004010040100401004010040100401004010040",
INIT_1A => X"FFBFBFFF7CFE7F9E79E7FFEDDFEFFFBEFFE7DF83F7EFFFFDF7E0000000000000",
INIT_1B => X"FDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FBFDFEFF7FB",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800003FFFFFF",
INIT_1E => X"8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8001000040000000000",
INIT_1F => X"FFFFFFFFFFD74AA552E80010552EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A",
INIT_20 => X"2ABDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A800105D2EBFFFFFFFFFFFFFFFF",
INIT_21 => X"FFBD54BA552A800100000001FFFFFFFFFFFFFFFFFFFFFFFBD54BA5D2E8201000",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF7FBD74BA5D2E800BA5D00001FFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A552A800BA5D2E821FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E820BA5500001FF",
INIT_24 => X"FFFFFFFFFEFF7FFD74BA552E801FF002E975FFFFFFFFFFFFFFFFFFEFF7FBD74A",
INIT_25 => X"00008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA552A8200014003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E80",
INIT_27 => X"BDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2E800005D2ABFFFFFFFFFFFFFFFFFF",
INIT_28 => X"BD54BA552E82028002AB8FFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2A80000412A",
INIT_29 => X"FFFFFFFFFFFFFFEFF7FBD74BA5D2A800281C00001FFFFFFFFFFFFFFFFFFFFF7F",
INIT_2A => X"52A820AA490A071FFFFFFFFFFFFFFFFFFEFF7FBD74AA5D2E800AA5500021FFFF",
INIT_2B => X"FFFFFDFEFF7FFD54BA5D2E80082492E871FFFFFFFFFFFFFFFFDFEFF7FFD74AA5",
INIT_2C => X"0000038FFFFFFFFFFFFFFFBFDFEFFFFFD54BA5D2A801C7142E955FFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8000008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005D043FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"54BA552A80010002ABDFFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2E800005D2EBF",
INIT_30 => X"FFFFFFFFFFDFEFF7FBD74AA552E820BA002AA8BFFFFFFFFFFFFFFFFFFFFF7FBD",
INIT_31 => X"E800BA5D04021FFFFFFFFFFFFFFBFDFEFF7FFD74AA5D2A800BA5504021FFFFFF",
INIT_32 => X"FBFDFEFFFFBD54BA5D2A820AA082A955FFFFFFFFFFFFFFBFDFEFFFFFD54BA552",
INIT_33 => X"52E975FFFFFFFFFEFF7FBFDFFFFFFBD74AA5D2E80000082A955FFFFFFFFFFFF7",
INIT_34 => X"00000000000000000000002ABFFFFFFFFFEFF7FBFFFFFF7FBD74BA552A801455",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"8632CA211E4491D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"24B000808800040439245B221373581F97B0A8D1040F92000F42000047A00E58",
INIT_05 => X"011B2BBA308F023810004700083E220811E9BF2844021B1004045E4249500449",
INIT_06 => X"80A51003AA0200C020088E16A85235722940A817251101010100040D6D0702A2",
INIT_07 => X"5C9ECAB0D247B013B405EAD525FAE48FC2060B880081A26DCD4047EFF9EF0189",
INIT_08 => X"2D0141C0055280100751096B6A40D6F86723E510AA2004803D3275EB2024E814",
INIT_09 => X"04804818CD280100207246A8020000AC0283002004051507A5411C0DA0005048",
INIT_0A => X"2C6898B2950AA65635B00041C23020131A80CFDFF3FE509A907C556828201102",
INIT_0B => X"050F60E220A06880D2A14050A028501428054278142151262CA50343854E506A",
INIT_0C => X"612B3482C0C0078E1F412B1582C090078E1F840A2B0114020104022460002200",
INIT_0D => X"012B1582C0C0078E1F412B3482C090078E1F891C239F8908003099C1ACF06273",
INIT_0E => X"1BA859F213AFC14AA380430060181BA1B0FD16770236A4091621C08055C2C0DB",
INIT_0F => X"B08AA600CA88B143AB11880C280600101F09C030AB28B03C111C239F87082804",
INIT_10 => X"4B61BD8068B92400D0004E30368910E8822A984B0025B0DE6089462660095337",
INIT_11 => X"001AC2173B00E162563454C40804055412D4481128C4CC012A66F30455309600",
INIT_12 => X"50840180A00E1C81900C4190E160589C48082C006A9057CA4385809520F07830",
INIT_13 => X"004416B105036B4180C000800C8C00460848952220592745AC11A544B1BF0068",
INIT_14 => X"512C6A8C4F0008AA800470370000A0004D0000002126F30C902A29C54539C020",
INIT_15 => X"2A81C2A81C2A81C2A81C9540E1540E001400006100003202D040050220103D2A",
INIT_16 => X"22365034A8EA754008004C0214202C50013456520CA09281C2A81C2A81C2A81C",
INIT_17 => X"104411044110441104411044110441104411044110441104411044110445E220",
INIT_18 => X"0401004010040100401004010040100401004411044110441104411044110441",
INIT_19 => X"0003FFFFFFFF9004010040100401004010040100401004010040100401004010",
INIT_1A => X"FFBFAFBEFDFFBBBEFBEFBEFBDFD1FE3EFBD7ADF9B3EFDF7DF7D0512289000000",
INIT_1B => X"FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79EFFC",
INIT_1C => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000FE7F3F",
INIT_1E => X"8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2A8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8201008043FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74AA552E80010552EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E8000055",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD54AA5D2A82000552ABFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2A800005D2EBDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A800105D2EBFFFF",
INIT_24 => X"FFFFFFFFFFFFFFBD54BA5D2E82010002AA8BFFFFFFFFFFFFFFFFFFFFFFFFD54A",
INIT_25 => X"0100004000000000000000000000000000000000000000000000001FFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001008043FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74AA552E800105D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A820001400",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD54AA5D2E800005D2ABFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A80000412AB8FFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A82010552EBDFFFFF",
INIT_2B => X"FFFFFFFFFFFFBD54BA552E80038492EB8FFFFFFFFFFFFFFFFFFFFFFFFBD54AA5",
INIT_2C => X"00000001FFFFFFFFFFFFFFFFFFFFF7FBD54BA552E82028002AA8BFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201000040000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74AA552A820005D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001000043F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD54AA552E8001055003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"A820105D2ABDFFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2E800005D2EBDFFFFFFF",
INIT_32 => X"FFFFFFFF7FBD54BA552A80010002AA8BFFFFFFFFFFFFFFFFFFFFF7FBD54BA5D2",
INIT_33 => X"02AAABFFFFFFFFFFFFFFFFFFEFF7FBD74BA552E800AA082EA8BFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000000021FFFFFFFFFFFFFFFFDFEFF7FBD74AA552E820BA0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"5886C0201A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"0005EE040057700F40D08078500000D9218020407F0000BB8018A2FC380BEAC2",
INIT_05 => X"FFE0419028700023FCBC385F87C0BFFFE0124002FFE1E0C517FF09111212F300",
INIT_06 => X"16D03FFC96102081020000020489019C430480241202080810FFDFE000000000",
INIT_07 => X"0001160A003475C8100123400E20E1F40F439647FF4807E189A477EF81DF0AF1",
INIT_08 => X"801008000007FEFFFB110140695812CC4188D58A0AAA10803448D0844FB71000",
INIT_09 => X"4201258112D4487FF8001010FFF7DE4000000003BFF8C25818080020017F0F94",
INIT_0A => X"0C024000004A9400000FFDFF50010103134CAFDF03BA18000F39900037C3EBFD",
INIT_0B => X"C02812F00429DC92C40002000100008000105400C00400100000A01800080100",
INIT_0C => X"A1CAF13F214001521001CBF03F21100152100801C17E61841950B1C10FFF57FF",
INIT_0D => X"01CBF03F214001521001CAF13F2110015210088528E00E02C8200A430A424202",
INIT_0E => X"02C86040902AC60BACDF0E02D02001C1C044006D0C94FB94320880603C420B80",
INIT_0F => X"00010AF5052419D196441902801430182800A018D9CA8000648528E00D124802",
INIT_10 => X"4D101808458A5602E000892029110445C19960A00026880C006739000009B003",
INIT_11 => X"1009408021144CB042F880100C0601844068880CE72000013600600332C14000",
INIT_12 => X"F80E02120018390320F050144CB241D0B9023402085020825132C8CB5B404030",
INIT_13 => X"C200400020224000405F7FFFE0008E17C0D240406519400500840A9524EE38A1",
INIT_14 => X"AC810033149249C433200180082A06FF907FC308181204800600000000001BFF",
INIT_15 => X"010C1010C1010C1010C10086080860840063090442A18001B188300C48907120",
INIT_16 => X"0100000000000004002403EFC10302219A41C1443243050C1010C1010C1010C1",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200010",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000080200802008020080200802008020080200802008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000000000",
INIT_1E => X"8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8001000043FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2A8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA552A8200000043FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A552A8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8201008043FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74AA552E8000055003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2A8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E800000800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA552A8001008043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52A8200014003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8200008043FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74AA552E820101C003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E800105D043FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000043F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2A8001008043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"A8200008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001000043FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74AA552A820005D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552",
INIT_33 => X"5003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA552E8200055043FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA552E800105",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"0000745C200801000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"0001E6000053300F00D0007810042140C00000407F0000BB800000DC3801EA00",
INIT_05 => X"FFE0000008700003FC3C380F87C019FFE01240009BE1E00003BF00000000F300",
INIT_06 => X"06103FFC000000000000000004890088010080001202000000FFDFE000000000",
INIT_07 => X"0009B24B043980021000810284204A8001401643FE4007E5501AA00000DC8C30",
INIT_08 => X"0000000000007EFFFB11A56940581280031D61420000B080102040BC5B006120",
INIT_09 => X"020125811254083FF80000003FF7DE0000000003BFF8005800000000017F0000",
INIT_0A => X"0000000000000000000FFDFF4000000AA0354000019C40000128000011C3EBFC",
INIT_0B => X"C000104000000010440000000000000000001000C00000000000000240058000",
INIT_0C => X"4012500021B00880108012500021E00880104809C1666594584031010FFF56FF",
INIT_0D => X"0012500021B00880108012500021E0088010492064206100E81084200048C080",
INIT_0E => X"0410004C840041A0D8005410903804100144800803419043064900C002050184",
INIT_0F => X"020902F60002260D65B361BAA1041018140F02C0000809408D20642053027004",
INIT_10 => X"00020818B06D9802F00030C02060110002C9E8010C00010480B35A0300400041",
INIT_11 => X"20042108603100061516EE800C060228204300166B4060080008240593D00218",
INIT_12 => X"7C02000040206602C10B48110006143B62023C00142800B04400095DFF902030",
INIT_13 => X"C000000000000000001F17FFE000DC1180C7804400044029208301040214AE4C",
INIT_14 => X"008000010012414433000100080806FD107FC300000000000600000000001BFF",
INIT_15 => X"000C1000C1000C1000C100060800608400630104408180012188300C00814080",
INIT_16 => X"0000000000000000000003EF80020201904181003003000C1000C1000C1000C1",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"F30C2416857732AEBAEBFFA55EDCF9822659AE7BE742E6441990000000000000",
INIT_1B => X"3C1E0F07BEFBEFBEF9E79E79E79E79E7BEFBEFBEFBEFBEFBE7BE7BE7BE7BEC98",
INIT_1C => X"83C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F078",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8000001E0F07",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008040000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8001000043FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2A8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008040000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2A8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008040000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8000008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000043FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8000008043FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A800100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00004000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"4909E6093253306F82D0007C80000000080E01007F8020BBC00040DC3801EA00",
INIT_05 => X"FFE0000008704503FE3C380F87C019FFF01241009BE1E00203BF80800000F392",
INIT_06 => X"06103FFF9E2086C2086E006604C9019D03108B741202605040FFDFE070400880",
INIT_07 => X"4024057000000100000000000000000001401643FE4007C00000000000CC0830",
INIT_08 => X"0801404000007EFFFF40010000401408000045000000A0801000408000000000",
INIT_09 => X"4A7DF795965C6D3FFC0020003FF7DF01880C618FBFFDD75E00100040437F0000",
INIT_0A => X"0000000000009400000FFDFFC006020000000000019804000028000191C3EBFF",
INIT_0B => X"C02812E0182000F2C48304418220C11160845004D04820000000000000000000",
INIT_0C => X"0002400001000800000002400001000800000801C0786184185031810FFF56FF",
INIT_0D => X"0002400001000800000002400001000800000000202000000800000000080080",
INIT_0E => X"0000000404000000880000001000000001000000000090000008000000040000",
INIT_0F => X"000100C600800001040000040009100000000200200000400000202000020000",
INIT_10 => X"0002000000081001000000000040010000082000000001000001080000000040",
INIT_11 => X"0080000040010000001080001008000000010000210000000008000010400000",
INIT_12 => X"0000030280000000010000010000001020000000000000100400000108000040",
INIT_13 => X"E0120012C1400080291F17FFF0018C11808200400000400000C2000000042000",
INIT_14 => X"00800001001243443B000100880806FD107FC301800000000600000000001BFF",
INIT_15 => X"000C1000C1000C1000C10006080060840077330C4889CC292588300C00804000",
INIT_16 => X"82068C0200000008014023EF80020201904189003003000C1000C1000C1000C1",
INIT_17 => X"110441104411044110441104411044110441104411044110441104451044C820",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FFFFFFFFFFFFC110441104411044110441104411044110441104411044110441",
INIT_1A => X"200A625D144BC2B4D34D7F61432D518B45265EF8278C2015DA080800002FFFFF",
INIT_1B => X"88C4623124924924924924924924924904104104104104104124904124904281",
INIT_1C => X"58AC562B158AC562B158AC562B158AC562B158AC562B158AC56231188C462311",
INIT_1D => X"00000000000000000000000000000000000003FFFFFFFFFFFFFF800002C562B1",
INIT_1E => X"8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"0003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"94A7B2B1450000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"6FEBEF5FEC737AFBC6F85FDEB220109E1FEFFFE3FBA7FDFB9BD301DC3FF5F0D2",
INIT_05 => X"FEEDBFDC387F987FEF7C3FAF87FF59F7F5FB7FF59BE1FF980BBBB7FE6D21F3DB",
INIT_06 => X"57902FFDEE9D7DC9D7DF2B263893479DDFAFDFE15213FEFEBFFFFBE1F1D3A333",
INIT_07 => X"10992310605CE10301DE0C1831CB7DF60A244B9BFEE00589DDBCEFEDC1DFA089",
INIT_08 => X"001D8EA111DA7FEFF90F21C8C84D9C0D858FC7020828C18FD18346BBF0000180",
INIT_09 => X"F37DF7B9DF7DCB3FDE89ECC07DF7DF5F985C6BCFFBFA28F99E7EB07F47FFEFAA",
INIT_0A => X"7DCFE1D4077B4D0026FFFFBE7D67D7F3BB79CFFB83BF14EC1E7D5980580BFAFF",
INIT_0B => X"C7D7D51D6F5FDCB935D7AFEBD7F5EBFBF7FEBD66DBFCA3F87501AE7B08060730",
INIT_0C => X"01F45EC0010007E01001F45EC0010007E010084BCD7FF1B61B5C33813FFFFCFF",
INIT_0D => X"01F45EC0010007E01001F45EC0010007E01001BD8020500008001F0100405202",
INIT_0E => X"1EC00040B02007EC09A0E00010001DC0004600400F781429C0080000770001A0",
INIT_0F => X"404B3BFD0402346235408402C08010003C064000E408010081BD802060020000",
INIT_10 => X"0E401A08FE0012040000FC002001360403E434588007200D00F88C84C081C203",
INIT_11 => X"001F01002156040675809145400007B00040091F1190982038406807C868B100",
INIT_12 => X"008320C0403C34000088601604067D00212000007C400082D81009FC08281D00",
INIT_13 => X"F7BFFED3FBFF6A84383F177FF005FFBFF5FA1040076065F730FC08043A903A80",
INIT_14 => X"F589807B7096CD4CF73AC1FC98884FFF19FFC71FEFED7B251E35768E8ED6BFDF",
INIT_15 => X"8C0D78C0D78C0D78C0D7A606BC606B8C56F7730ECCDBDF152199F51EDDCDEBCF",
INIT_16 => X"DFE7DD87FEFF7FF796FFFFFDFFD7E681B867D3683A03A40F78C0D78C0D78C0D7",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFEFDFD",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"FFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEB",
INIT_1A => X"57AA9ABAD8ACBF0E38E3A89F9E923C2CD990A7D0D2A377F86EDB5C88646FFFFF",
INIT_1B => X"4C261309861861861861861861861861861861861861861861A69A6986186EBC",
INIT_1C => X"84C26130984C26130984C26130984C26130984C26130984C26130984C2613098",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000261309",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"1085B0B041000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"6FAB975B6470BAF386C87A9CB00000001FEF9F23E3A7BDE79B5101D23FB5C0C2",
INIT_05 => X"F8EDBFD4347F18778E723F2E47FE59C7F5FB7F759B91FB880BA3B6FE2921CBDB",
INIT_06 => X"47000FFC128D5CE8D5CC210638A046889CAB57E8421786B6ACFFE3E181932377",
INIT_07 => X"000000042000000288020C18300320620A80231BFE200181092CE7ED80DFC001",
INIT_08 => X"000C562551D87E8FF90041101042110180004102800008801183468180000141",
INIT_09 => X"137FF7A0FF75813F1C85244071EFBF17D85C738BE3FA08F9DE36B05B07FEEF22",
INIT_0A => X"768EA0C406630D00226FFE3E2D62D6E21259CFDB039E806C02451880400BE0FC",
INIT_0B => X"CC57550D63564D1D2556ADAB56D5AB6AD7EAB962CBD8A3A83101F47E08040510",
INIT_0C => X"01E44A40010007600005E44A4001000760000843C561E5C55C42B9011FFF48FF",
INIT_0D => X"05E44A40010007600005E44A40010007600004BD8020100008001F0100001302",
INIT_0E => X"1EC00000382006EC0820A00010001DC0000208400D781020C008000077000020",
INIT_0F => X"40431BC50402146235400400408010003C064000C400018080BD802020020000",
INIT_10 => X"0E400204FE0010040000FC0000003E0403A424108007200102E888808081C200",
INIT_11 => X"001F0100005E040475808101400007B00000015D111010203840081748482100",
INIT_12 => X"00012040403C34000080201E04047D00202000007C400000F81001FC08080500",
INIT_13 => X"E5ADA4C25ADE72041A3F147FF0018DBBB5FA10400360649310FC08003A903A80",
INIT_14 => X"054880693016DD4C755AC16C1A884FFE18FFD757E7ED7A211E81C09818109E1F",
INIT_15 => X"440C3440C3440C3440C3C2061A2061AD46FF730E5CCBCD55219AB55F0DEFABC7",
INIT_16 => X"5EC71385FC2512E3565BBBF1BAD6F281BC63F1683803C00E3440C3440C3440C3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BDE75ED",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"FFFFFFFFFFFFAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB",
INIT_1A => X"200E5E48710A4200000028150200903950C086D0E28028104A471688747FFFFF",
INIT_1B => X"0080402000000000000000000000000000000000000000020800000000000780",
INIT_1C => X"5028140A05028140A05028140A05028140A05028140A05028140201008040201",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8000028140A0",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"8C2100804900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"02000100440408002408008002221000204116A280000F000001400000100010",
INIT_05 => X"0004D44400004D4400000000000000000000005C0000000A0000002C20600000",
INIT_06 => X"4100000120040A0040A00B0090006202940100004000A2020400200888800911",
INIT_07 => X"5002489020420110800244891211440804000810002000081040000000200000",
INIT_08 => X"080542C004CA00000050080202008401842004108AAAA00008912240A1248804",
INIT_09 => X"0000000C0000E400002040500000009202C1002040004400022200020400B062",
INIT_0A => X"58C460540329810002D002000400407020800000004000640800088008280001",
INIT_0B => X"0140000401028008330000800040002002480102010082981500062108020430",
INIT_0C => X"00040A40000000A00000040A40000000A0000040060084104110828030000800",
INIT_0D => X"00040A40000000A00000040A40000000A0000000800010000000000000005000",
INIT_0E => X"00000000A00000040020A000000000000006000000080020C000000000000120",
INIT_0F => X"4040152000000020000004004080000000000000240000000000800020000000",
INIT_10 => X"0000120002000004000000000001220000040410800000090000808080800002",
INIT_11 => X"0000000001420000200001014000000000000900101010200000480008082100",
INIT_12 => X"0001204000000000000820020000200000200000000000028800002000080500",
INIT_13 => X"00933050080C0001900020000000408010000000022000D61028000008000000",
INIT_14 => X"400082D022040000400800081022C0000080000206CB0821082B694D4D294000",
INIT_15 => X"050160501605016050160280B0280B0012000843066021001400040024440245",
INIT_16 => X"0861CD33548542A10209D4100E4040A00002002C004001036050160501605016",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008021081084",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"0000000000000020080200802008020080200802008020080200802008020080",
INIT_1A => X"06A0A0F108816B1861863BED822140048D2E5818732C5589A40A0C22E1000000",
INIT_1B => X"80C0603020820820820820820820820820820820820820820820820820820035",
INIT_1C => X"582C160B0582C160B0582C160B0582C160B0582C160B0582C16030180C060301",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800002C160B0",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0803B2814D0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"26E1E905CC574828C4F85FC600000016004F77E2F887CDB80BC340DC07D1F000",
INIT_05 => X"FE1DFE4C080F884FE33C078F803F19F011E93ED49BE01F1A03B8972E6D20F049",
INIT_06 => X"57902000DE142D4142D5030010134395D70589415002DA4A17FFF800F0C38111",
INIT_07 => X"00092300601CE00101DE040811D919F402244293FEE00400CCB46BA4C164A088",
INIT_08 => X"08148A4000887FE0000F20C8C80D080D818FC2000000418FD08142BAD0000884",
INIT_09 => X"E204D2154D28AA3FC60888D03C10415A80402847F8002458926A002E457FA0AA",
INIT_0A => X"5587A1540231410006DFFF80540541619968C76980E914E4163D4980100BFA02",
INIT_0B => X"07C7C0140D0B50A8218102C0816040B1225C1506512C83E85500AC3A08040630",
INIT_0C => X"00141EC0000000A01000141EC0000000A01008480D3EB4A24A0C910037FFFC00",
INIT_0D => X"00141EC0000000A01000141EC0000000A0100100800050000000000000405200",
INIT_0E => X"00000040B000010401A0E000000000000046000002080429C0000000000001A0",
INIT_0F => X"40483B590000202000008402C080000000000000240801000100800060000000",
INIT_10 => X"00001A08020002040000000020013600004414588000000D00108484C0800003",
INIT_11 => X"000000002156000220001145400000000040090210909820000068008828B100",
INIT_12 => X"008320C00000000000086016000220000120000000000082D800082000281D00",
INIT_13 => X"32936E43A92F2880B01F37001004B29450580000066021F6303C000408000000",
INIT_14 => X"B481806A62840800C22800B8900042FF0180000ABFEF89250815568A8AD6ABC0",
INIT_15 => X"8D0068D0068D0068D006A68034680300021410028450530014014002D445624D",
INIT_16 => X"89418D13FE7F3FFD8BADB7FC4F4164A00806522C0A40A50268D0068D0068D006",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C4B12C9894",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"FFFFFFFFFFFFC0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0",
INIT_1A => X"FFBF3F5E7CFC7DFFFFFFD7FADDCFFFBEFFCF1F879DFFFFFDFFEA0C00602FFFFF",
INIT_1B => X"DFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBAEBAEBAEBAEBAFFFD",
INIT_1C => X"FDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800003EFF7FB",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"F7AEBEBFFDFFBFBEFBEFFFFFDFF3FC3EFFF7FDFBF76FF7FDFFD0000000000000",
INIT_1B => X"FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79EEBD",
INIT_1C => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000FE7F3F",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"1084B030000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"6DA986092050306382C05A1C900000001FAE89016387B2A38B5000D03FA1C0C2",
INIT_05 => X"F8F92B90307F41338E303F0E07FE19C7F1FB7F289B81FB8003A396D20940C3DB",
INIT_06 => X"06000FFC020004C0004C000628800488080003600213001000FFC3E101030222",
INIT_07 => X"000000000000000220000810200220620E00030BFE000181092CE7ED80DF8001",
INIT_08 => X"0000000001107E8FF90001000040100000004102200000801102448100000100",
INIT_09 => X"027DF780DF74013F1C00240071E79F05888C618BA3F800599C101049037E4F40",
INIT_0A => X"240A808004420400202FFC3E002202021259CFDB039E0008024510000023E0FC",
INIT_0B => X"C407500020004C10060204010200810040801060C04821202001A05A00040100",
INIT_0C => X"01E04000010007400001E0400001000740000803C0616184184031010FFF40FF",
INIT_0D => X"01E04000010007400001E04000010007400000BD0020000008001F0100000202",
INIT_0E => X"1EC00000102006E80800000010001DC0000000400D7010000008000077000000",
INIT_0F => X"000308C50402144235400000000010003C064000C000010080BD002000020000",
INIT_10 => X"0E400000FC0010000000FC000000140403A020000007200000E808000001C200",
INIT_11 => X"001F01000014040455808000000007B00000001D010000003840000740400000",
INIT_12 => X"00000000403C34000080001404045D00200000007C400000501001DC08000000",
INIT_13 => X"E004048240426200081F147FF0018C1380DA10400140640100D4080032903A80",
INIT_14 => X"050800A91012494C31004124080886FE187FC301B124F2001600000000001A1F",
INIT_15 => X"000C1000C1000C1000C18006080060840477330C4889CC012188310E08812982",
INIT_16 => X"02061004A820104809402BE1900222019861D1403803800C1000C1000C1000C1",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100446020",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"FFFFFFFFFFFF8100401004010040100401004010040100401004010040100401",
INIT_1A => X"00000000000000000000000000000000000000000000000000001000802FFFFF",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000000000",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"88280C4C7B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"00160090920C04800904848262220277E05152B280780D407428E723C01E1400",
INIT_05 => X"0006D46207801E400183C0707800E6000E008057641E00473C40680D32330C00",
INIT_06 => X"C165000225E2C11E2C12A0D0144AC27206582C166504816162002000B0FC21D5",
INIT_07 => X"5E6D233B964E7CD99DFB870E1DDDD889C5FBDC440129A0604442180238203F70",
INIT_08 => X"AD23C17544C581000657A0E8E83D86F0E4A7B2D88AAAFD7FE0E1833AC5920CFC",
INIT_09 => X"6D82082E2081B6C0027ADA398000008A504318404005B70663212C04A080B036",
INIT_0A => X"414568729139FA5610C00001A2502440888420247041E87681008CE9AFC80001",
INIT_0B => X"22B826E250B12346F1244812240912048941621804A150CA1CA45C254D4AF4AA",
INIT_0C => X"F80FA97FE0F0009E0FC40FA97FE0F0009E0FC048211E9C11C31F82E4A0008900",
INIT_0D => X"040FAB3FE0F0009E0FC40FAB3FE0F0009E0FCC42EFDFBF0AE03080E2AEB2E0F1",
INIT_0E => X"013879BA878FE807F65FBF12E0380231F0BD9E3FC08FEBD6F661C0E008C3CB5F",
INIT_0F => X"B248831ACBFC8BBDCAB779BC699F20180309A0F83BE2B87C7C42EFDFBF187806",
INIT_10 => X"4131B59003FFEC07F00003F01FB90BE9F01FC8B38C2098DAE007F323A0C83136",
INIT_11 => X"3080E29F1B2BE9F8A27E6E915C0E004C72BEC800FE7464290626D7003F994718",
INIT_12 => X"FC0C2352A0024B83F07F198BE9F8A0FFDA2A3C0202B8776A2FA7F023F7D06570",
INIT_13 => X"1448126105810941C5C068000CD4004C0905E52630BB1AE49C2BA7F98D6F846D",
INIT_14 => X"6074EA560F0416A24844B01302A26100C4801844069B0C88881A28C141118000",
INIT_15 => X"A781E2781EA781E2781C33C0613C0E21020800239450116ED443C041B47E9665",
INIT_16 => X"241140A056954AB0C280D0002020187007122C3E04E03383E2781EA781E2781E",
INIT_17 => X"20481204812048120481204812048120481204812048120481204812058112C1",
INIT_18 => X"0481204812048120481204812048120481204812048120481204812048120481",
INIT_19 => X"0000000000001204812048120481204812048120481204812048120481204812",
INIT_1A => X"C4109CAF9C4C83B8E38E2AE9C136AD8E9B562CF042E6281CF13043A85D400000",
INIT_1B => X"F0F87C3E08208208208208208208208208208208208208208208208208208220",
INIT_1C => X"1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1",
INIT_1D => X"000000000000000000000000000000000000C3007FFFFFFFFFFFA00000F87C3E",
INIT_1E => X"4214555517DEAA5D7BFFEAAF7803FEBAF7FFD74BAAAAABDEBAF7AE8000000000",
INIT_1F => X"1555FF55517FE000055421FF00557DF45A2D5401EFF7D142145A2AE800BA0851",
INIT_20 => X"5555555A2AABFFFF5D516AA00A28028A00AAAEBFE00A2FBD75FFFF8400155085",
INIT_21 => X"5517FF45A2AEBDEBAAAAAA8BFFF7D140010FF84174BA552EBDFFF0004020005D",
INIT_22 => X"5504000BA5D2E97545A28028B4508554014508043FEBA082ABFE10AAAEA8ABA5",
INIT_23 => X"FA2AABFE00FFFFD74AA085540000002E801FF557FD75FF0051401FF5D0015410",
INIT_24 => X"EFF7FFC20BAF7D1575450800020BA08517FF45F7FBFFF45A2FFFDE00002E801F",
INIT_25 => X"A38BF8FC000000000000000000000000000000000000000000002ABEFAA80001",
INIT_26 => X"7155BC2A87092AAFA9257F1C5BC00AA5D7FF8EAA57803AEBAF7F5D74AAA2A03A",
INIT_27 => X"BFBC7EB8005B55A85B555EF095F50578085BE8FC7A3F00516DA2D5451D7EBDB4",
INIT_28 => X"0975FFAAA1521FF492BF8F40B6AAB84AF555168A00EA8000150A801C01C7142E",
INIT_29 => X"2EBAE28168ABAA2D43D568BC5400168E90E2F412BEAE3D542A004380124921D2",
INIT_2A => X"2FA3AA28EA8168A954100071D2E90A855C7A00A38F6DE05B40480557A95A3A1C",
INIT_2B => X"16D1EAE925EA0BFEBF4AA09217F490568417085147B50A80095178157FEFA074",
INIT_2C => X"000002D57AAA8402A8743DBD202DA95568A95E800A8F57F6DA971F8F7FFFA42D",
INIT_2D => X"AAFFD1564BA2282BFA02A2C28000000000000000000000000000000000000000",
INIT_2E => X"5EFA87F57555AAFBD7555FFAE95408A8FDC31AD017D34ABA5D7BEAAAAD786BCE",
INIT_2F => X"C2087383F79A5046A37B55F38415555797D63BFF007F8B2B2D97D483AFA7BD9F",
INIT_30 => X"42000D382964A92B401E71D7581C33172EC0A0300A6AEA8FAF0451CA001D4845",
INIT_31 => X"C8365A2FD5E04AA5780A8AAAD7AC3CA02003BEBBA7D7463CC508D07577BAFBD5",
INIT_32 => X"0621F562B1122DA70C3808458881056A5502AA150502828811FCD4EABDB1DFDF",
INIT_33 => X"96D55BBAAC55EAFAF86D35E4A92B4460D15060374FF72AAADF24559515705079",
INIT_34 => X"007FC0000007FC0000007FC07AAF12E00505D3FDF6A03D4BFB79AFA4C5CB5F58",
INIT_35 => X"0007FC0000007FC0000007FC0000007FC0000007FC0000007FC0000007FC0000",
INIT_36 => X"00000000000000000000000000000000000000007FC0000007FC0000007FC000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000040000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"CA1800080848B0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000010822C00803804000001999EF9C00040B0002000001000640200001018",
INIT_05 => X"0000400244000000014200004000000004000000001000032000200002100800",
INIT_06 => X"208500000080412804100CB08000302220080408010000202000000404100844",
INIT_07 => X"5AF6FEF002230018010860C1833C460044204C000008A0041000080008202800",
INIT_08 => X"8D22C0F55000010000524481890BC000263000188AAAA10F8C1830562B25FC4C",
INIT_09 => X"B102002E20013600022D8819000000A000110A4000002C204000240420001000",
INIT_0A => X"02605C1C1108481200C000002040040820000020104100028800002801041001",
INIT_0B => X"081001004010810510040802040102008100200800A1100707040101E20BE0B0",
INIT_0C => X"58000003C0F000A000C4000003C0F000A000C0000012187087010AE4B0000000",
INIT_0D => X"04000003C0F000A000C4000003C0F000A000CC4200002F08E03080000010F180",
INIT_0E => X"0000000AAC00680000001F10E038000000078808C00000023461C0E000000127",
INIT_0F => X"5200040A00D000000202090C281F201803000000240218C0044200001E187806",
INIT_10 => X"400012900001EC03F000000000392100B00048230C200009A000130320480002",
INIT_11 => X"308000000961002880204A901C0E00000002C9000260640900004D0000904618",
INIT_12 => X"5C0C0312A002000000083881002880025A0A3C020000002A8400B00007806070",
INIT_13 => X"04080830008010468220A00008D0000801046004308A18500002012800090428",
INIT_14 => X"0840280206089000004090110200000000001454000200828008081110084000",
INIT_15 => X"4191AC191AC191A4191A00C8560C8D2910000060901010401E13405111220000",
INIT_16 => X"0410028000100800140000002004103224002006406401918C191AC191A4191A",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200800041",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"0000000000000200802008020080200802008020080200802008020080200802",
INIT_1A => X"2431A589945201924924B060D757DF8A94102E038728287452B4008A04000000",
INIT_1B => X"75BADD6EAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8A28A28A28A28AB20",
INIT_1C => X"974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D6EB75BADD6EB",
INIT_1D => X"00000000000000000000000000000000000303FFFFFFFFFFFFFFC00000BA5D2E",
INIT_1E => X"FDFFFA2FFD74000855555FFFFFFC01FF087BE8BFF5D2AAAB5555554000000000",
INIT_1F => X"EBFF455D04175FF5D7FEAAAA002ABDEAA5D2EBFFEFA2D17DEBAF7D1574BAAAFB",
INIT_20 => X"8415400005540155F7D16AB45002EA8ABA005540145557BFDEAA5500154AAAAA",
INIT_21 => X"5003DE00A2FFFFFEFAAD57DE00082AAAA00082A820BAAAD540145F7D5574BAAA",
INIT_22 => X"F7D5554AA5D2ABDEBA082A821455D2EA8B455D2A975EFF7AEBFF550055555FF5",
INIT_23 => X"FFF84155FFFFFFFFF55AAAABFFFF5D556AB45A2D16AABAAAAEBFE10AAFBD7545",
INIT_24 => X"10FF84174BA552EBDEBA0004020AA5D04155FFAAFFEABEFA2FBEAB455D7BD55F",
INIT_25 => X"F47015A800000000000000000000000000000000000000000000175FFF7D1400",
INIT_26 => X"FEAAF7D5524AAA2F0BAF7FABDFC7E10005F525D74BFBC51FF1471E8BEF55242F",
INIT_27 => X"50492490E17EAAA2AAB8F4515043DFC75575C7000B6AEBAEAA5D2EBDFFFBED17",
INIT_28 => X"B6FB6DF7DFD5038ABA140A2D00554517DEBDB6FB55142A8708202FBD257F1C75",
INIT_29 => X"AABFF55BC5B555C74B8A38E38085BE8B47A3A00503D1420AD000B420820AAE2D",
INIT_2A => X"AABD21EF1C2FEA5FDEBDB505FA4920AFE10082E925555F8FFDE38087FC51C7F7",
INIT_2B => X"1EFBFDBFF5FF1C00BF5D25475C7B7FEAFF45BEAABA4AF555168B68FEDF6AB52A",
INIT_2C => X"00000151EAE3D542A004380124921D20BFFFA0AA17AEB8BFF155552B6F5E8BFF",
INIT_2D => X"FF55516ABEFDD003EFE5093DC000000000000000000000000000000000000000",
INIT_2E => X"2BA5D2ABDFFFF7D57DEAAFFD5420B2A2D37DB07A3D795000087BC01458AFBC11",
INIT_2F => X"D608897FD610D01151C610592A974BAFBAC28B55550434D555C53E0CE2AAA874",
INIT_30 => X"3FE102400144ABAAFFF7DE772FDD56588042F72EF0851575FFAAFBDD5542B2ED",
INIT_31 => X"F6A81A239501755F504BDF557D79431FD006EABA100F3D68FFFAABAC20EF0400",
INIT_32 => X"55EAF57FF957CAAA7FABF7DFD0C6A7DFFFA07FC04EA0006BFE007E2E8315DD02",
INIT_33 => X"FADF6900FFFF68BEFDFFB4B1FE5551141E78A02803158517BD745AEAEA8FAF0C",
INIT_34 => X"0000000000000000000000165BAFBD542000D382964A92B403EE18D5408A6F2A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000040000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0812",
INIT_01 => X"A145A00810790848048044A54E404340404000720885800802000906E4910200",
INIT_02 => X"5C010802020408040C455850AA055254090541A111200A104A0000000908B510",
INIT_03 => X"182002200C00004485264A001214912802150020218808002440854288890550",
INIT_04 => X"210302008014100120806B08702010102722C9E0412200651102418214049492",
INIT_05 => X"48416A98042912208552102442884882A58A08011290A1120A81230240018DCA",
INIT_06 => X"12800554528021C8023A28000031240048000100001170000155414109102066",
INIT_07 => X"000022104040810089080810211A04480420420154800088096A0EA8C0222080",
INIT_08 => X"080198C105424705510A08828A0B19080428040080A0A10F8102049300000804",
INIT_09 => X"3165541CD54822160A89E89020AA8AC4CA1D39CE215264B04040002400B80688",
INIT_0A => X"280201840548C80001C568146000001012D40D7182411080153801004800B057",
INIT_0B => X"4812050000080114100206000100818100900640C04C20104101021C00000310",
INIT_0C => X"00A00000010000A01001400000010000A0100801407234E34C1A980001552055",
INIT_0D => X"01400000010000A01000A00000010000A0100038000000000800000000405000",
INIT_0E => X"00000040A00002600000000010000000004608000850000000080000000001A0",
INIT_0F => X"400020C4000200420040000000001000000000002408000000A1000000020000",
INIT_10 => X"00001A04940000000000000020012800018000000000000D0288000000000003",
INIT_11 => X"0000000021480000508000000000000000400951000000000000681300000000",
INIT_12 => X"00000000000000000008600800004C000000000000000082A000015000000000",
INIT_13 => X"80004012C06000018004342AA000700000000000044000500000000022101800",
INIT_14 => X"958100134200904487400010022005E0110D524029263100009200151409130A",
INIT_15 => X"C9013C9011C90134901144801A4808AD4451394CD0391A541593C04B59084008",
INIT_16 => X"010400A0A890684444240120C0071420344423040240450114901149013C9011",
INIT_17 => X"080601806018060180200802008020080601806018060180200802048026C000",
INIT_18 => X"8000080001804018040180400800008000080601806018060180200802008020",
INIT_19 => X"1F83F03F03F00180401804018040080000800008000180401804018040080000",
INIT_1A => X"E90C042CB002102CB2CB2EE00271AE180616A85246C77250C7D00022012F81F8",
INIT_1B => X"28944A2504104104104104104104104104104104104104104104104104104608",
INIT_1C => X"128944A25128944A25128944A25128944A25128944A25128944A25128944A251",
INIT_1D => X"000000000000000000000000000000000003C3007FFFFFFFFFFFCE3F00944A25",
INIT_1E => X"EAA1055042AA105555421EFFFD568AAA002EBFEBA550002000AA800000000000",
INIT_1F => X"AA8BEFAAAE975FFA2D5555450851574000851554BAFFAE801FF087BE8BFF5D7B",
INIT_20 => X"2EA8AAA5D2EBFFFFA2D1554BAF7D17FEBAAAFFFDFFFA2D57DE10557BE8ABAF7A",
INIT_21 => X"D04175FFFFD5574AAAAAA974BA082EA8BEFAAD555555F7D568ABAF7D5574BA55",
INIT_22 => X"085557410F7AA97410087BD55FF087FEAA10A2FFEAAAA552AAAAAAAAAABFF455",
INIT_23 => X"05D7FE8B45F7FBFDE00085540155F7D56AA00007FEAA000055401555D7BFFE10",
INIT_24 => X"00082A820BAAAD540145F7D557410AA8428A10550017400550402155A2803FE0",
INIT_25 => X"000E28A80000000000000000000000000000000000000000000017400082AAAA",
INIT_26 => X"01FF1471E8BEF5574AFA00010ABFA38555F401D74BD16FAAA002ABFEAA550E82",
INIT_27 => X"FF400417FEF082F7AAA8BEFE2AA955EFA2DB5757FEAFBD2410005F57482E3AA8",
INIT_28 => X"F6DA82F7DF520385D2FE80AA5D2EBDFD7BED1574AAF7D5524AAA2F1FAF7FABFB",
INIT_29 => X"24ADAAAB6AAB8F455784155C75575C7000B6AE95492082EADBFFBEDB55555E3D",
INIT_2A => X"051C05571474024A81C5557578EBA087400007FC21C7005B6FB47F7A438E925D",
INIT_2B => X"E10A001FFB40038F68F7F578F7FFEF568E2808554717DEBDB6FA3D0075EDA800",
INIT_2C => X"000001043D1420AD000B420820AAE2DB4716DF7DFFDE381D716FA15550015428",
INIT_2D => X"AA002ABDEAA552A80010AAA88000000000000000000000000000000000000000",
INIT_2E => X"800087BD5410AAAA801FF55556ABEF5D517EEE00828FDEBA5D7BC015582D57DE",
INIT_2F => X"A2B2A3D169B07A3D7BFE10597BFDE00AEAC28BFFAAAE955EFAAFBC15F5A3D7D6",
INIT_30 => X"BDFEFFFFBC1154AAFFFFE107FF9D72A20842080BA5D2ABDF55F7D575EAAFFD50",
INIT_31 => X"97CF4780286A2105D2A3FEBAFFAC28B555504145555A53C00B2A2AA02000082A",
INIT_32 => X"FFFDA02003FFDEAA8557D65550915544AA5D51574EAA28015400547FC315D007",
INIT_33 => X"16F9E2555500174AA282E20BFFFF842AAAAADD5699ADABD5A8AAA0051575FFA2",
INIT_34 => X"0000000000000000000000030EF04003FE102400144ABAAFFD75E7F2BDDD2B80",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000080000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380202",
INIT_01 => X"200C9A424080216D3C2462C99E104B49404040028804A0080A000416A8D90A0C",
INIT_02 => X"4809A902031800444461089C66E331352180D468B8240E600C0081110B80ACD0",
INIT_03 => X"DA16C2210C0001D231A30A0648C68428320066010A80881068A80C401CC46330",
INIT_04 => X"2088601DA82700EC92307064A3756910088469A01C250210990240420E005A48",
INIT_05 => X"2D2060182414411A314A0A02C18C01B9854368080A506912018C2502484038D1",
INIT_06 => X"16801CCCAA8061E8061C0D008020140520080769000420202133CCC50C110804",
INIT_07 => X"5800B65040630008810C20508138071604A461833280038C89904E6400232008",
INIT_08 => X"0800906010521D1CC80204918949540C061000088000A90F840A50963A017845",
INIT_09 => X"A037A02C68552A35620C88900A69876100810A6A84C82C400040300D40D20A48",
INIT_0A => X"062A10B40042C80000CCE4CC2045051913208CE80243048008204100402079CC",
INIT_0B => X"C81301004C18912102060C0207010201C190200400A401042D00F15884030170",
INIT_0C => X"0190148000000800100450148000000800100401CB33494594532980733322CC",
INIT_0D => X"05101480000008001004F014800000080010051C000040000000000000480000",
INIT_0E => X"00000044000001680180400000000000014000000B1004090000000000040080",
INIT_0F => X"00812E44000024400140800280000000000002000008000001B0000040000000",
INIT_10 => X"0002080CCC0002000000000020401000034010480000010402D8040440000041",
INIT_11 => X"00000000601000064180104400000000004100570080880000082015C0209000",
INIT_12 => X"00820080000000000100401000061C0001000000000000904000094C00201800",
INIT_13 => X"4408400000A26285A03224E670094008010000004444010E2050000420801880",
INIT_14 => X"4DC10283429294408740C0B48202854C011CD75C0102A30400A8891451284B26",
INIT_15 => X"4901A4901849018C901A648056480C2D4449116DC0115C41159B655F112AC008",
INIT_16 => X"0510000000DA690C1D20030BA0011421B404220402404501A49018490184901A",
INIT_17 => X"280803808038080380803808038080380C0280C0280C0280C0280C0680C28051",
INIT_18 => X"00C0280E030080380A030080380A030080380C0280C0280C0280C0280C0280C0",
INIT_19 => X"B556AA9556AA830080380A030080380A030080380A0200C0280E0200C0280E02",
INIT_1A => X"742C000A981E80249249206018F18E0C85142822266800586291000A844D54AA",
INIT_1B => X"A9D4EA7524924924924924924924924924924924924924904104104104104A20",
INIT_1C => X"1A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A753A9D4EA753",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF849010D46A35",
INIT_1E => X"42000AA802AA10F7D57FEAA557BE8B45A2D5555EFAA800015508000000000000",
INIT_1F => X"BC0155A280021EFA2FFE8B4555042AA105555421EFFFD568AAA002EBFEBA5551",
INIT_20 => X"D5574000851554AAFFAE801FF087BC01FF5D7FEAA10550402000AAD56AAAA557",
INIT_21 => X"AAE975FF005540145A2D157410AAD17DFFF5D0400010AA842AAAAFFD542000FF",
INIT_22 => X"F7AE975FF080428B455D7FFDEAA5D55574BA00517DE105551420BAF7AAA8BEFA",
INIT_23 => X"F007FFFEAAAAD5554AA552EBFFFFA2D5554BAF7803DEBAAAFFFDFEFAAD57DEAA",
INIT_24 => X"EFAAD555555F7D568ABAF7D5574BA552E800BAAAAE800AA087BD5555552A821E",
INIT_25 => X"155080E800000000000000000000000000000000000000000000020BA082EA8B",
INIT_26 => X"FAAA002ABFEAA555E02000E28AA8A38EBD578E82E975EAB6DBEDF575FFAA8E02",
INIT_27 => X"87A38AAD56DA824975C217DAA84021FFAAF5EAB55EBAEADA38555F451D7EBD16",
INIT_28 => X"E2DABAFFDB47412ABFE90410005F57482E3AA801FF1471E8BEF5575EFA00012A",
INIT_29 => X"5F47082E3AAA8BEFA02A955EFA2DB5757FEAFBD2400BED57FFD7410E05038BE8",
INIT_2A => X"2F1FAF7FABFBEAE2AEBA4974871C043AB6D4975FFEBA5D71D742A407FFFE0055",
INIT_2B => X"1C75D25C74920821D708757AE2AA3FFC04AA552EBFFD7BED157482F7803AEAAA",
INIT_2C => X"0000007092082EADBFFBEDB55555E3DF6DA82F7DF7AE38497FC00BAB6A485082",
INIT_2D => X"FFFFFFD75FFAAAE8014500288000000000000000000000000000000000000000",
INIT_2E => X"EBA5D7BD5545A2D57DEAA002EBDEAA557BC0010AAA8A8ABAAAD568A1020516AB",
INIT_2F => X"29EF5C517EEE00828D74AAFBD57DE000057C21FFAA80001FFAAD57EB55A2A8AB",
INIT_30 => X"7DF55082E974AAFFAABDEBA77FDD66A0ABBDC2000087BD5410AAAA801FF55556",
INIT_31 => X"7C14100957FF6105D7BD5400AAAC28BFFAAAE955EFA8FBC15E5A3D5D7400FFD5",
INIT_32 => X"D1554A8FFC42AA10A7D169F57ABD7FEEBAAA841550555002ABFF54517EEB25D5",
INIT_33 => X"96F014AAFF84154105555C215500000014558557FA42A3D7020BA5D2ABDF55F7",
INIT_34 => X"000000000000000000000015400082ABDFEFFFFBC1154AAFFFFE10FFF9DF2020",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000040000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204002",
INIT_01 => X"010398000008004C1C20650E1E104348403008418984014902030006A0910200",
INIT_02 => X"480108A200000000444048E41E80F00A4104311868200200080000000988A390",
INIT_03 => X"0CA08220080000D004060A0240101028270012603000000030808C0208C000F0",
INIT_04 => X"4403A609A055306BC2C0735810CEE5100A0A40E06B8360E3808241D03845D002",
INIT_05 => X"ECE0498800791403AD3038AE079059A790E245819A41E4120BAB87800001D312",
INIT_06 => X"06000C3D220003E0001A210088B1008C4004034912120000010FC3C00000A064",
INIT_07 => X"5000220440000000090800002118400204206100F040018019004B8001232088",
INIT_08 => X"0810884441123323C0424180880B0108002000000880890F9000041200000845",
INIT_09 => X"230B6715A4786E0F5A8C889031EF9F45D884794FA03A24781840100D000E1140",
INIT_0A => X"0C4202200142400004DC3C82600401003200872003FB1400082840001022003C",
INIT_0B => X"C800940008088034040000010000808140901000C00001008800A01814000840",
INIT_0C => X"02E0100000000800000620100000000800000001C07261841840310240F070C3",
INIT_0D => X"0680100000000800000760100000000800000435100040000000000000080000",
INIT_0E => X"00000004000000D8008000000000000001000000155000080000000000040000",
INIT_0F => X"000100EC00004002214000008000000000000200000000000094100040000000",
INIT_10 => X"000200010C000200000000000040080005800008000001000368000040000040",
INIT_11 => X"000000004008000448000040000000000001007C000008000008001D00001000",
INIT_12 => X"000000800000000001000008000017000100000000000010200002C800000800",
INIT_13 => X"0000549000027200800E271E00288400800208004804C0080000000052800800",
INIT_14 => X"454000924280D144B14041340A880EC51160525C0022510006BE1002C6150F5E",
INIT_15 => X"010C1010C1010C3010C14086980861AD447F2201D899BA403593514B59A30088",
INIT_16 => X"010448002098694C15204369E00116203445E3443043410C5010C3010C1010C3",
INIT_17 => X"180000006018000000200804010020080400002018040000600800010064E000",
INIT_18 => X"8060000001000008060180201000000040180001006008000100201804000020",
INIT_19 => X"934D964C32698000401802008060000401000008060080201004000000080201",
INIT_1A => X"0991A185145019A28A289830C700FC0A0002870BB5ED0B34504048828464B261",
INIT_1B => X"351A8D46AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8A28A28A28A28AF4C",
INIT_1C => X"8341A0D068341A0D068341A0D068341A0D068341A0D068341A0D46A351A8D46A",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8EE3EC1A0D06",
INIT_1E => X"40155080000155FF843FFEFAA84001FF5D043FEAA5D55420AA002A8000000000",
INIT_1F => X"A80010FFAE975FFAA80001EFA2AAAAA10F7D57FEAA557BE8B45A2D5555EFAAD1",
INIT_20 => X"AAAAA105555421EFFFD568AAA002EBFEBA555542000AA80001555D04174AA002",
INIT_21 => X"280021EFA2FFE8B45F78400145FF842AAAAA2AA800BA5D51555EF002AA8BFFAA",
INIT_22 => X"00003DFEF080428B455D002AABA5D2AAAAAA5D2E82000AAD568AAA557BC0155A",
INIT_23 => X"FAAAAA8BEF552E820000851554AAFFAA801FF087BC01FF5D7FEAA105D0428B45",
INIT_24 => X"FF5D0400010AA842AAAAFFD542000FFD57DF55A280154BAA2FBE8AAAF7AA821E",
INIT_25 => X"092142E00000000000000000000000000000000000000000000015410AAD17DF",
INIT_26 => X"AB6DBEDF575FFAADE02155080E85145E3803FFEFA284051D755003DE92415F42",
INIT_27 => X"851455D0A124BA002080010FFA4955C7BE8E021C71C0A28A38EBD57DE824975E",
INIT_28 => X"B505D71424AABD7F68E2FA38555F451D7EBD16FAAA002ABFEAA555F42000E2AA",
INIT_29 => X"D56DA824975C217DAA84021FFAAF5EAB55EBAE82145F7802AABAA2A480092415",
INIT_2A => X"575EFA00012ABFB6D080A3AFEF080A2FB45490E2AA824924AAA92550A07038BE",
INIT_2B => X"AAFFEAA00F7AE821D7B6A02FBC71D0E10010005F55482E3AA801FF1471C01EF5",
INIT_2C => X"0000010400BED57FFD7410E05038BE8E2DABAFFDB6FA12ABAEBDF7DAA80104BA",
INIT_2D => X"4555043FE10087BC2000552C8000000000000000000000000000000000000000",
INIT_2E => X"ABAAAD57DE1000516ABFFFFFBD75FFAAFFC0145002897555A2803FFFFAA84175",
INIT_2F => X"DEAA557BC0010AAA895555042E820BA080400010FF8017545F7AE821455D2CAA",
INIT_30 => X"2AAAAAA8002010007FC0155D5022A955FFACBFEBA5D7BD5545A2D57DEAA002EB",
INIT_31 => X"43CAB0552C97CAAFFD57DE000057C21FFAA80001FFAAD57EB55A2A880155F780",
INIT_32 => X"AA801FF5555421EF58517EAB00028A9BEF002EAABEF002EBDF45542AAAA00080",
INIT_33 => X"A90FDFEFA280020BAA2FFEAA10FFAE82145F7803CFE55D2CC2000087BD5410AA",
INIT_34 => X"000000000000000000000002000FFD57DF55082E974AAFFAABDEBAF7FDDE6A0A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000080000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A337A20E07C0C1E006",
INIT_01 => X"295FBC448000804C5C6A60000C34C26841280A00084000C8C212802EE2953235",
INIT_02 => X"C809AD5EB118E640A4D158FC011FF0002080000082E8C66609DB7DDDCB1FA036",
INIT_03 => X"4A120E4C3A4C90D214A35E824852857A0A20640A88800000B8E0FC52A884500E",
INIT_04 => X"001440809A2604005934800041110A71E290E8B010DB221C662AE22DC0AA3448",
INIT_05 => X"12026A2A1B88C31841CDC451B860A6507BEBD18A65AE10571450DE8112522449",
INIT_06 => X"80752C03736281D628398CD0A4C894EA2054237F271331095100D82D0C2C82A2",
INIT_07 => X"5E64B66BD6231CC81529A356AD3AC601C57FF54FF149A46490261C4B39203F70",
INIT_08 => X"AD0099410015814FC602C4B1B93947F8621030C800001D7FA46A95172E937835",
INIT_09 => X"2C836D35B68D26C082DE9AB88C104020000208401807B78739010C04E17F5014",
INIT_0A => X"082099129008F25615C3FC01A2102109204C28B6706168128920C469E7C00A00",
INIT_0B => X"E92C23E210A0B246C2234010A108D0042811461C0401502644A40106C14FD22A",
INIT_0C => X"E00BF1BFE1F000BE1FC40BF1BFE1F000BE1FC80028120800800100653FF0313F",
INIT_0D => X"040BF53FE1F000BE1FC40BF53FE1F000BE1FCC806FFFEF0AE83080E2AEF2F1F1",
INIT_0E => X"013879FAAF8FC003FEDF5F12F0380231F0FF963F00A7FBDF3669C0E008C3CBFF",
INIT_0F => X"F2008022CBAC8B9DDEB779BEA91F30180309A0F83FEAB8FC7C006FFFDF1A7806",
INIT_10 => X"4131BF940DFFFE03F00003F03FB929E9C19BE8EB0C2098DFE2EF7B2760483137",
INIT_11 => X"3080E29F3B69E9F4427EEED41C0E004C72FEC95DEFE46C090626FF1537F15618",
INIT_12 => X"FC0E0392A0024B83F07F7989E9F01DFFFB0A3C0202B877EAA7A7C1CBFFD07870",
INIT_13 => X"C0404020040001C4E7F1787E0C8028514885C566241902508C83A7D1B7EFAC6D",
INIT_14 => X"4DF46A170F92C7E20F0430938008AC38C4184B100136858C9298A8560688F4C1",
INIT_15 => X"6B8C86B8CE6B8CA6B8CC15C6435C670C10EB4124D2B3903BF5C9710C1191DCA0",
INIT_16 => X"2030461200984D041C40208400230E71B3104E5636E3178C86B8CC6B8CA6B8CE",
INIT_17 => X"0040118401184610042110401184410846110421104010844118421504238200",
INIT_18 => X"8441184011844100461004211046100461084211042100441084011842100461",
INIT_19 => X"DA6924965B4D1004610840118401084410840110421004610046110421084410",
INIT_1A => X"FF9FBFAF2DDA3B9E79E7BED9CFEF73B6FFE74FC3F78FFF6DB7ED438A183124B2",
INIT_1B => X"DDEEF77BBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEDFD",
INIT_1C => X"BDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BB",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF853FB5EEF77B",
INIT_1E => X"020AA002AAAABA555140155087FFFFEF00042AB555D2E955FFF7FFC000000000",
INIT_1F => X"E975FF5D5568B555D7BD5545FFD540155FF843FFEFAA84001FF5D043FEAA5D04",
INIT_20 => X"FFEAA10F7D57FEAA557BE8B45A2D5555EFAAD5401550800001FF5D00001555D2",
INIT_21 => X"FAE975FFAA80001EF002AAAABAF7D168A10A2D17FF45A2FFC0000AAAE974AAFF",
INIT_22 => X"F7803DF55FFAEBFE005D2EAAB45557BD55555555401555D04174AA002A80010F",
INIT_23 => X"5552E955EF5D7FEAA105555421EFFFD568AAA002EBFEBA555542000A28028BFF",
INIT_24 => X"AAA2AA800BA5D51555EF002AA8BFFAAAA820AA5D517DF55082E974BA087FE8B5",
INIT_25 => X"5C7F7FBC0000000000000000000000000000000000000000000000145FF842AA",
INIT_26 => X"51D755003DE92410F42092142E28ABA5D5B4516D007FFFFFF1C042FB7D492A95",
INIT_27 => X"851C75D0E02145492E955C75D5F6DB55497BD5545E3DB45145E3803AFEFA2840",
INIT_28 => X"BC7028A2AA95492FFFFE8A38EBD57DE824975EAB6DBEDF575FFAADF42155082E",
INIT_29 => X"0A124BA002080010FFA4955C7BE8E021C71C0A2DABAF7D16DA28A2DB7AF7DB6F",
INIT_2A => X"55F42000E2AAA8BEFE3843AF55E3AABFE105520AFB45557BD5555415F4514549",
INIT_2B => X"082E954AA087FEDB7D5D2A155D7157BEFA38555F451D7EBD16FAAA002ABFEAA5",
INIT_2C => X"0000002145F7802AABAA2A480092415B505D71424821D7F68E07082495B7FF7D",
INIT_2D => X"EF5D003DFEF002E95555F7FDC000000000000000000000000000000000000000",
INIT_2E => X"555A2802ABFFAA841754555043FE10082A82000552CAAAAA5D7FD75EF087BFDF",
INIT_2F => X"75FFAAFFC0145002895545552E80145002E955455D7BFDF45007FD7555A2F9D5",
INIT_30 => X"7FEAAAAFFEABFFF7FFD54BAA2AA95410F7FDEAABAAAD57DE1000516ABFFFFFBD",
INIT_31 => X"BD55550879D5555002E820BA080400010FF8017545F7AE821455D2CBFEAAFFD1",
INIT_32 => X"D57DEAA002EBDEAA557BC0000AAA8A8BEFA28028B45AAAABFE0009043FF555D7",
INIT_33 => X"FAC97400087FFFFFF002E954AA087BFFFFF5D2E975455D7DFFEBA5D7BD5545A2",
INIT_34 => X"000000000000000000000000155F7802AAAAAA8002010007FC0155550222955F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000300000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B0061A258A2840112C03002C180004003220200403302301C0381A0082",
INIT_01 => X"860041C838394848008100000042026041000000090800090210010000510204",
INIT_02 => X"080108220C1000004464080000C008010000000001243240080080000988A050",
INIT_03 => X"080000010C23404080020A600200002983800504488000103080050C08C10000",
INIT_04 => X"0040504280A682104011230010000010002040E9102050101000400A00003000",
INIT_05 => X"0409400984008000414A00014000002004100020005004020010204044802800",
INIT_06 => X"301223FC028911E8911900000224200248A653E908C0248489FF000809108000",
INIT_07 => X"0000220441820000090C080001184400142040200E824008900008000220600A",
INIT_08 => X"1A18946451007FA0380200808809010C182000000000090F8100001220000804",
INIT_09 => X"300240B4A409223F020988100808200490142B441BF82C20401481540A000008",
INIT_0A => X"264285180542408000D001BE090693912000002004410489080001100017E2FD",
INIT_0B => X"091081090A4491A40052A129519428CA142288010A5A21214601F01A220602A0",
INIT_0C => X"18100400000000A00034100400000000A00033A00813004104020818800F2400",
INIT_0D => X"F4100080000000A00034100080000000A0003142000000000000000000055D00",
INIT_0E => X"00000001E8002900010000000000000000066000C20004000000000000000120",
INIT_0F => X"4D240C2000502000000080000000000000000000240146800142000000000000",
INIT_10 => X"00001260F0000000000000000007F00032201000000000091A00040000000002",
INIT_11 => X"0000000005D00008958010000000000000003F4000008000000048D240008000",
INIT_12 => X"008000000000000000082670000CC0000000000000000007C000301400200000",
INIT_13 => X"0120849A5250101482202301F05101202420000810C219500150002800101280",
INIT_14 => X"454110030212C140011204D020880C000018431DE802015022A62A1596C8B580",
INIT_15 => X"016C2016C2016C6016C440B6000B600C446B0104D09192013589701C59800002",
INIT_16 => X"51804A0028904C425016040820978221B0000005B05B416C0016C0016C4016C4",
INIT_17 => X"8CA3294A528CA328CA1294A528CA3284A5294A728CA3284A529CA728CA100508",
INIT_18 => X"CA3284A129CA7294A328CA1294A729CA128CA329CA5294A128CA3294A5294A32",
INIT_19 => X"1C71C718638E28CA529CA7284A128CA7294A528CA1284A729CA1284A3284A529",
INIT_1A => X"ED9DBDAFBC5E9BBEFBEFBEF9CFF1FE1E9F52AFF9F3E77B7CF7F40A00107638C3",
INIT_1B => X"FCFE7F3F8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E76C",
INIT_1C => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9",
INIT_1D => X"00000000000000000000000000000000000303007FFFFFFFFFFFC61AC8FE7F3F",
INIT_1E => X"955FFF7FFC21EFF7D17DEAA5D2AAAAAA5D557DE105D2EBDF55557FC000000000",
INIT_1F => X"03DEAA5D5568BEF5D042AA10A2AAAAABA555140155087FFFFEF00042AB555D2E",
INIT_20 => X"5540155FF843FFEFAA84001FF5D043FEAA5D00020AA002A82145555542010FF8",
INIT_21 => X"D5568B555D7BD5545FFD568AAA5D00154AAAAD1420BA00557DF455D7BFFEAA55",
INIT_22 => X"F7843FF55007FFDEAAA284020BAAAD168BFF0800001FF5D00001555D2E975FF5",
INIT_23 => X"5AAAEBFE10FFFFEAA10F7D57FEAA557BE8B45A2D5555EFAAD540155080000000",
INIT_24 => X"10A2D17FF45A2FFC0000AAAE974AAFFFFC21EF5551401EFF7842AA00FF841754",
INIT_25 => X"F45497FC000000000000000000000000000000000000000000002AABAF7D168A",
INIT_26 => X"FFFF1C042FB7D492A955C7F7FBC71EFFFD57FE825520ADA92495B7AE10412EBF",
INIT_27 => X"0716D415F47000F78A3DE92415F6ABD7490A28A10AAAAA8ABA5D5B4516D007FF",
INIT_28 => X"F78F7D497FFFE925D5B45145E3803AFEFA284051D755003DE92410E02092140E",
INIT_29 => X"0E02145492E955C75D5F6DB55497BD5545E3DB6AA92550A104AABED1470AA005",
INIT_2A => X"ADF42155082E87038FF8038F6D1C7BF8EAAAA80020BAA2DB68BC7140E051C75D",
INIT_2B => X"FF8428A00E38412545AAAE3FE10A3FBE8A38EBD57DE824975EAB6DBEDF575FFA",
INIT_2C => X"000002DABAF7D16DA28A2DB7AF7DB6FBC7028A2AA95492FFFFC71EF415F471C7",
INIT_2D => X"00007FEAA10002ABFF450079C000000000000000000000000000000000000000",
INIT_2E => X"AAA5D7FD75EF087BFDFEF5D003DFEF002E95555F7FDD55EFF7D57DE005D003DE",
INIT_2F => X"FE10082A82000552C955FF007BD5410FFAABFE00087BE8B45082EAAA10A2A8AA",
INIT_30 => X"820AAF7D5574AA087BEABEF007FFDE00557DD5555A2802ABFFAA841754555043",
INIT_31 => X"BEAB55552C95545552E80145002E955455D7BFDF45007FD7555A2F9EAA005D2A",
INIT_32 => X"516ABFFFFFBD75FFAAFFC01450028974BAFF842ABFF557BE8ABAA284020BAA2F",
INIT_33 => X"7FDD55EF007BD5555F7802AA10AA8000145AAAEBFE10A2F9EAABAAAD57DE1000",
INIT_34 => X"00000000000000000000003FEAAFFD17FEAAAAFFEABFFF7FFD54BAA2AA95410F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000240000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C024504188000003000000003302300C018180006",
INIT_01 => X"020008422008604D042080000211024840000000080000080200080000110204",
INIT_02 => X"4801082048100000444008040080000041000000000222400800000009000010",
INIT_03 => X"0802030288A148D0000208424000002103006400088000003080000408C10000",
INIT_04 => X"00004000890600004032030010000010008060E4100000140006500800403040",
INIT_05 => X"0400400080000018414800810000002000000000004000328010000080882000",
INIT_06 => X"281A8001220021E0021803000224200200000360888420000000100808000000",
INIT_07 => X"5000220409020000090800000118040014A061200052500810000C490323208E",
INIT_08 => X"1A9098411110014000424090980B0002102000000000010F8000001220000805",
INIT_09 => X"31024034A4092200820D899408000004D0143B4410002C800080020450800001",
INIT_0A => X"24028011444240A88CC00100200D0010200008B2066397014800221400140C01",
INIT_0B => X"080001000C008124000000000100008000100404204C25200451A01A00A620A5",
INIT_0C => X"1C0014800000F001E02C0014800000F001E021141213000000000010B0001000",
INIT_0D => X"CC0014800000F001E02C0014800000F001E022420000400004C3201C51040908",
INIT_0E => X"60078601084038000180400002C0E00E0E004100E000040900000B0380383400",
INIT_0F => X"08146800105100000000800284004160C0301D07001504820242000040000198",
INIT_10 => X"908C404AFC000200030F000FC00610103BE0104810C8462014F8040446120C88",
INIT_11 => X"C3201C608410100FD5801044013098038D00309F008088C2419100A7C0209021",
INIT_12 => X"00B2048902C0807C0E008450100FDD000100411C8107880440403DDC00201804",
INIT_13 => X"00100496406010A0A2002200125140000000221110C018066250402E32901A80",
INIT_14 => X"454214028220141530400910CA800900326790500002001444001C0050140A00",
INIT_15 => X"5120551205512055120708901A8901A104804000801212541403C15178008010",
INIT_16 => X"01004200A09A49445420000DC000152804C9A384814809201512015120151201",
INIT_17 => X"0004000000080200806008020000000000000020080200802000000000008000",
INIT_18 => X"0000000000802008000000000002008020000400000000000080600802008000",
INIT_19 => X"0002082080000100000802008020100000000008020180000000000020180200",
INIT_1A => X"0000000000000000000000000000000000000000000000000005428A14584104",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8DD9EC000000",
INIT_1E => X"BDF55557FFDE00557BEAABAA2AEAABEFF78015555AA801741055554000000000",
INIT_1F => X"BEAAAAAAD157555AA803FEBA5555421EFF7D17DEAA5D2AAAAAA5D557DE105D2E",
INIT_20 => X"802AABA555140155087FFFFEF00042AB555D2E955FFF7FFD5555557BEABFFF7F",
INIT_21 => X"D5568BEF5D042AA10A2AA955EFF7FFD5400F7FFFDFEFAA80000BAAAAA820BAA2",
INIT_22 => X"5D7FE8A000004154BAF780001EFAAAAA8B45000002145555542010FF803DEAA5",
INIT_23 => X"5AAD5555EF557FC0155FF843FFEFAA84001FF5D043FEAA5D00020AA002ABDEBA",
INIT_24 => X"AAAAD1420BA00557DF455D7BFFEAA5555575455D2AAABFF5551421FFAAD15754",
INIT_25 => X"4385D5540000000000000000000000000000000000000000000028AAA5D00154",
INIT_26 => X"DA92495B7AE10412EBFF45497FFFE385D71E8AAAAAA0A8BC7EB8417555AA8410",
INIT_27 => X"D056D5D75EABC7FFF5EAAAABEDF5257DAA8438EBA4155471EFFFD57FE825520A",
INIT_28 => X"0070BAA2A0870BAAA8028ABA5D5B4516D007FFFFFF1C042FB7D492A955C7F7FB",
INIT_29 => X"5F47000F78A3DE92415F6ABD7490A28A10AAAA925EFEBFFD2400EBFBFAFEFAA8",
INIT_2A => X"10E02092140E3DE924171E8A281C0E10482F784001D7AAA0AFB6D1C040716D41",
INIT_2B => X"4955421EFA2DF5557DAAD5D05EF0175C5145E3803AFEFA284051D755003DE924",
INIT_2C => X"000002AA92550A104AABED1470AA005F78F7D497FFFE925D5B525454124AFBC7",
INIT_2D => X"55A28015545A284000BA5D534000000000000000000000000000000000000000",
INIT_2E => X"5EFF7D57DE005D003DE00007FEAA10002ABFF450079FFEAA5D5568ABAA2842AB",
INIT_2F => X"DFEF002E95555F7FDC01EF55556AB55F7D56AABAF7FBC01EFA2842AABA085755",
INIT_30 => X"C2000A2FFEABFFAA84174BAAA80174AAAA862AAAA5D7FD75EF087BFDFEF5D003",
INIT_31 => X"43DFEF5D02155FF007BD5410FFAABFE00087BE8B45082EAAA10A2A8801FFA2FF",
INIT_32 => X"841754555043FE10082A82000552CBFE10085168AAA552A80010F78000145AA8",
INIT_33 => X"57DC014500003FF450051401FFA2FBD55EFAAD5421FF085755555A2802ABFFAA",
INIT_34 => X"00000000000000000000002AA005D2A820AAF7D5574AA087BEABEF007FFDE005",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0000040042840002C00000018000002700500030B3132000400812082",
INIT_01 => X"A14008420008204D042100000212026840000000180800080200090048510200",
INIT_02 => X"080108020090000004655C000080000051000000002402400800000009008010",
INIT_03 => X"0002000100300C408422420002108108028065044880001030808D4288C10000",
INIT_04 => X"0002504688A28210003100000000001002A0E88910A032541000090A00643040",
INIT_05 => X"04092A081400D118410A002140004020140001A9005000004810A1C0044D2800",
INIT_06 => X"0010EFFD228931C8931820002080258A48A653E00213248C98FFC0094910A222",
INIT_07 => X"4000220440120000090C0810210A040034A040000046180810000C4907036008",
INIT_08 => X"50D88C2450000140004200808809000C012000000000010F8102041320000000",
INIT_09 => X"2002002020010200828C88020800200040801A40100228A1585481544A804040",
INIT_0A => X"A20804802400C80080D0010029069290200008B20E2304086800400640200801",
INIT_0B => X"091084090A4C81240251A328D094684B34A288050A5828012009504420102180",
INIT_0C => X"080004801E0FF00010000004801E0FF000100220021200000000000080001000",
INIT_0D => X"000004801E0FF00010000004801E0FF000100440000000F517CF600000400104",
INIT_0E => X"E000004008100800010040ED0FC7E000004008804000040109963F1F80000080",
INIT_0F => X"0020040020100000000882431660CFE7C0F00000000800810040000000E587F9",
INIT_10 => X"B0000808000001F80FFF0000200008021040134473D800040010045C1F360001",
INIT_11 => X"CF600000200802028001102EA3F1F80000400002008B83D6C0002000802688E7",
INIT_12 => X"03F2DC2D1FC18000000040080202800004D5C3FD80000080200818000027928F",
INIT_13 => X"0122C01A52501094222002000110012064200008848218002100100C00004112",
INIT_14 => X"4500048240C08400841204D0A00089000100001DE9248104300294428148A480",
INIT_15 => X"4800048000480004800004002240020850884000901210140011C010312B888A",
INIT_16 => X"51A4C000889A4D0E1D7624086491800420044240020004004480004800048000",
INIT_17 => X"84A1284A128CA328CA328CA328CA328CA328CA1284A1284A1284A12C4A14E508",
INIT_18 => X"CA328CA3284A1284A1284A1284A328CA328CA328CA328CA3284A1284A1284A12",
INIT_19 => X"000000000000284A128CA328CA328CA328CA3284A1284A1284A1284A328CA328",
INIT_1A => X"4799B1A014503EB65B6594F14A87D78AF421448BB528AF75D640088884400000",
INIT_1B => X"7C3E1F0F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79EDFC",
INIT_1C => X"87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F0F87C3E1F0F8",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF834FA53E1F4F",
INIT_1E => X"174105555420000000021EFAA843DE00F7803FEBAFFFFC2000557FC000000000",
INIT_1F => X"43DE005504175FF08514014555557DE00557BEAABAA2AEAABEFF78015555AA80",
INIT_20 => X"7FC21EFF7D17DEAA5D2AAAAAA5D557DE105D2EBDF55557FD54AAA2AA955FF000",
INIT_21 => X"AD157555AA803FEBA55556ABFFA280154BAFF803DF45FFD17DFFFFFD56AA0055",
INIT_22 => X"002AAAAAAA2D57DF450004154BA087BEAAAAF7D555555557BEABFFF7FBEAAAAA",
INIT_23 => X"5FFD1555EFA2802AABA555140155087FFFFEF00042AB555D2E955FFF7FFD5410",
INIT_24 => X"00F7FFFDFEFAA80000BAAAAA820BAA280000AAA2843DE1008556AA00A28028B5",
INIT_25 => X"0285D75C00000000000000000000000000000000000000000000155EFF7FFD54",
INIT_26 => X"8BC7EB8417555AA84104385D5542038000A001C7A2803AE38FF843DEBAEBFFC2",
INIT_27 => X"D24BAA2AA955C708003FE285D00155FF0055451555D5F7FE385D71E8AAAAAA0A",
INIT_28 => X"B78FFFE3DF6DA284175C71EFFFD57FE825520ADA92495B7AE10412EBFF45497F",
INIT_29 => X"75EABC7FFF5EAAAABEDF5257DAA8438EBA415568BEFA28E124AAF7843AF7DEBD",
INIT_2A => X"92A955C7F7FBD54380020ADA82BED57DF450804104920875EAA82F7DB5056D5D",
INIT_2B => X"005F68A10BE802DB55E3DB555FFF68028ABA5D5B4516D007FFFFFF1C042FB7D4",
INIT_2C => X"00000125EFEBFFD2400EBFBFAFEFAA80070BAA2A0870BAAA80070BAA2803DE00",
INIT_2D => X"AAFF803DEBAAAFBC20BA55514000000000000000000000000000000000000000",
INIT_2E => X"EAA5D5568ABAA2842AB55A28015545A284000BA5D53420BA082E82155AA802AA",
INIT_2F => X"AA10002ABFF450079C20BAAAAE9754500043DEBA5D04175EF0855575455D7BFF",
INIT_30 => X"820AAFF802ABEFAAFFEABEFAAFFFDEAA0051555EFF7D57DE005D003DE00007FE",
INIT_31 => X"16AA10FFFFC01EF55556AB55F7D56AABAF7FBC01EFA2842AABA085768BFFA2AE",
INIT_32 => X"7BFDFEF5D003DFEF002E95555F7FDD74BA08043DE10F7D17FF55000000010085",
INIT_33 => X"A86174AAAA843DE00087FE8A00F7843FF45AAFFD75EFF7842AAAA5D7FD75EF08",
INIT_34 => X"0000000000000000000000001FFA2FFC2000A2FFEABFFAA84174BAAA80174AAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000100000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000006",
INIT_01 => X"000009801830084C182060000C104268413C0A61590001D90213C00000110200",
INIT_02 => X"680108200010000054400C000080000041000000010002400800800009082011",
INIT_03 => X"0008000004002040000200100000000042800584488000103081880008800000",
INIT_04 => X"00005842802AC210001000000800001000004080100040140080040800003100",
INIT_05 => X"0400000040000080410800010001002000000000004000002010000040002000",
INIT_06 => X"10100001221911E1911902000020200201A2D3E8000C2C84880010080800004C",
INIT_07 => X"C0002204000200000B080000010C040004A0400000C0000810000C5901036000",
INIT_08 => X"002A84300000014000C2008088090000002000000000030F8000001220000408",
INIT_09 => X"210000020000120082088801080020400000084010002880000C803400000008",
INIT_0A => X"020000040000480100D0010019019190200008B2022380800802010000000801",
INIT_0B => X"09000119064C810500D0A36851B428DA14368C801A1400000100500400000090",
INIT_0C => X"08100080000000A00000100080000000A00000000212000000000000B0001000",
INIT_0D => X"00100400000000A00000100400000000A0000540000000000000000000005100",
INIT_0E => X"00000000A8000900000040000000000000060000420000010000000000000120",
INIT_0F => X"4000040000102000000000020000000000000000240000800140000000000000",
INIT_10 => X"00001204FC000000000000000001280013A000400000000900E8000400000002",
INIT_11 => X"0000000001480004D5800004000000000000091D008000000000480740200000",
INIT_12 => X"0002000000000000000820080004DD000000000000000002A00011DC00001000",
INIT_13 => X"0322C01032301006022082000010032024200000048019500000000832901A80",
INIT_14 => X"4501000200089400007200D0020008000000144C4800000200BC228404020080",
INIT_15 => X"0010000104001000010440080000822900000000801010500A13404111008000",
INIT_16 => X"D1A0CA0000984D06403600086591900224002000400440104001040010000104",
INIT_17 => X"8DA368DA3685A1685A1685A1685A1685A1685A1685A1685A1685A1685A120D08",
INIT_18 => X"5A1685A1685A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA36",
INIT_19 => X"000000000000685A168DA368DA368DA368DA368DA368DA368DA368DA1685A168",
INIT_1A => X"6C20080AB9A28724904120E1999E91BCD151200802001038E2550A0010100000",
INIT_1B => X"68341A0D14514514514514514514514514514514514514534D34D34D34D344A1",
INIT_1C => X"268341A0D069349A0D069349A0D068341A4D268341A4D268341A0D068341A0D0",
INIT_1D => X"00000000000000000000000000000000000003FFFFFFFFFFFFFF8A6AC8341A4D",
INIT_1E => X"C2000557FEABEFA2D1400AA5D2AAAA00F7FFEAA10F7D17FFFFAAAE8000000000",
INIT_1F => X"03DFEFF7FFE8ABAF7802ABEFAAAE820000000021EFAA843DE00F7803FEBAFFFF",
INIT_20 => X"843DE00557BEAABAA2AEAABEFF78015555AA80174105555421EFF78028BEF5D0",
INIT_21 => X"504175FF0851401455555555EFA2FBC01FFF7AAAAB45557BC0155007FFDEBAAA",
INIT_22 => X"552A974AAA2843DEAA5D2A820BA000428AAAAA84154AAA2AA955FF00043DE005",
INIT_23 => X"AF7D1400BAAAAE821EFF7D17DEAA5D2AAAAAA5D557DE105D2EBDF55557FFDE00",
INIT_24 => X"BAFF803DF45FFD17DFFFFFD56AA00557FC201000517FFEFAAAEBDF45FFAEA8AB",
INIT_25 => X"FD7A2A48000000000000000000000000000000000000000000002ABFFA280154",
INIT_26 => X"AE38FF843DEBAEBFFC20285D75EFBC7A2DB400824120ADA38E3F1EFA28F7DF7D",
INIT_27 => X"421C7FF8028BEF41003FFD7F7F1EDA82F78E2DBD7A2A482038000A001C7A2803",
INIT_28 => X"1C716D1475FFEAAA28E3FE385D71E8AAAAAA0A8BC7EB8417555AA84104385D55",
INIT_29 => X"AA955C708003FE285D00155FF0055451555D5F575C7A2FBC51EFEBA0A8B6D557",
INIT_2A => X"12EBFF45497FFFE105D2E97482AA8038EAA412E850AA1C0428ABAB68E124BAA2",
INIT_2B => X"B6A0BFF55F7AEAAA82FFDF40092B6A4871EFFFD57FE825520ADA92495B7AE104",
INIT_2C => X"0000028BEFA28E124AAF7843AF7DEBDB78FFFE3DF6DA284175C001000557FFEF",
INIT_2D => X"AAA2D57FEAAF7FBFDF45AA800000000000000000000000000000000000000000",
INIT_2E => X"0BA082E82155AA802AAAAFF803DEBAAAFBC20BA55517DF55A2FBC201008003DE",
INIT_2F => X"5545A284000BA5D5340145F78028BFF08003DF45FFD57FE00FFAABFF45AA8002",
INIT_30 => X"D75FFA2842ABFF5555575FF55557FEAAA2AABFEAA5D5568ABAA2842AB55A2801",
INIT_31 => X"028ABAF7AA820BAAAAE9754500043DEBA5D04175EF0855575455D7BD5555A2FB",
INIT_32 => X"003DE00007FEAA10002ABFF450079FFE005D2A97400A2802AABA002A954AA5D0",
INIT_33 => X"0514200008517DFEFFF803FF45FFAAA8A00F7FBC2010FF80155EFF7D57DE005D",
INIT_34 => X"000000000000000000000028BFFA2AE820AAFF802ABEFAAFFEABEFAAFFFDEAA0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000200000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110204",
INIT_02 => X"0801080200100000046558040080000041000000002402400800000009008010",
INIT_03 => X"00020201040000D0842242024210810802006400088000003080054288C10000",
INIT_04 => X"0000400088020000003020002000001002A0E881108032100002000800203040",
INIT_05 => X"04092A081000411841480001000000201000012800400010001081C040402000",
INIT_06 => X"10100001220001E0001802002020240208000369001520080100100909000266",
INIT_07 => X"4000220440020000090C0810210A040004A0410000C0000810000C4901036008",
INIT_08 => X"0000802100100140004200808809000C002000000000010F8102041320000000",
INIT_09 => X"2000000000000200828888800808000410800840100220211850004442004048",
INIT_0A => X"240A80800442400004C0010000060210200008B2022304880800410000200801",
INIT_0B => X"0000010008008020020100008000400120800004004821202001A05A00040180",
INIT_0C => X"08101400000000A01004101400000000A0100000081300410402080080003000",
INIT_0D => X"04101080000000A01004101080000000A0100540000040000000000000405100",
INIT_0E => X"00000040A80009000180000000000000004608004200040800000000000001A0",
INIT_0F => X"4000282000102000000080008000000000000000240800800140000040000000",
INIT_10 => X"00001A00000002000000000020013000100010080000000D0000040040000003",
INIT_11 => X"0000000021500000800010400000000000400900000088000000680000009000",
INIT_12 => X"008000800000000000086010000080000100000000000082C000100000200800",
INIT_13 => X"040004924040008020000200101100004000000000C019500050000800000000",
INIT_14 => X"4541008240801000804000108280800001001051A12481041080801010000080",
INIT_15 => X"4800048004480044800044000240022100884000901210440003C141102B088A",
INIT_16 => X"00044280009048485D4020080000140004046240020044000480044800448000",
INIT_17 => X"080200802008020080200802008020080200802008020080200802048026E011",
INIT_18 => X"0000000000000000000000000002008020080200802008020080200802008020",
INIT_19 => X"0000000000000080200000000000000000000000000000000000000000000000",
INIT_1A => X"CA83332A34488A8A28A29E195281FC1A72E24C2BF5A4D9555204428290100000",
INIT_1B => X"94CA65328A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A354",
INIT_1C => X"994CA6532995CAE572B94CA6532994CA6572B95CAE532994CA6532994CA65329",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF838CF1CAE532",
INIT_1E => X"7FFFFAAAE801FF08557DF4555516AA00007BEABEFAAD1555FFF7840000000000",
INIT_1F => X"56AA0000043FFEFA2FFFDE1008556ABEFA2D1400AA5D2AAAA00F7FFEAA10F7D1",
INIT_20 => X"84020000000021EFAA843DE00F7803FEBAFFFFC2000557FC0010AAD57FF45A2D",
INIT_21 => X"7FFE8ABAF7802ABEFAAAEA8BFF5D0415400F7FBFDEAA007FEAB45AAAE800AAF7",
INIT_22 => X"5D0415555557BFDFEF00517DE00A28028B450855421EFF78028BEF5D003DFEFF",
INIT_23 => X"A5D7FFDEBAF7AEBDE00557BEAABAA2AEAABEFF78015555AA80174105555401FF",
INIT_24 => X"FFF7AAAAB45557BC0155007FFDEBAAA8417410AAFFD7555AAD56AB45A2AE800A",
INIT_25 => X"5C7E380000000000000000000000000000000000000000000000155EFA2FBC01",
INIT_26 => X"DA38E3F1EFA28F7DF7DFD7A2A4801EF085F7AF6D55556AA381C75EABEFBED157",
INIT_27 => X"C0010AADF7AF6DB6D56FA3814003AFFFA2F1F8E381C516FBC7A2DB400824120A",
INIT_28 => X"5E8B45BEA0850BAE38002038000A001C7A2803AE38FF843DEBAEBFFC20285D75",
INIT_29 => X"8028BEF41003FFD7F7F1EDA82F78E2DBD7A2A4ADBEF550412428F7F5FDE92087",
INIT_2A => X"A84104385D55401C75504125455575FAFD7145578E10AA802FB450851421C7FF",
INIT_2B => X"BED56FB45BEA082082557BF8EBAF7AABFE385D71E8AAAAAA0A8BC7EB8417555A",
INIT_2C => X"00000175C7A2FBC51EFEBA0A8B6D5571C716D1475FFEAAA28E10438AAF5D2545",
INIT_2D => X"BA5D5568BEFF7D157555AA800000000000000000000000000000000000000000",
INIT_2E => X"F55A2FBC201008003DEAAA2D57FEAAF7FBFDF45AA80021FF007BE8BFF5D516AA",
INIT_2F => X"DEBAAAFBC20BA555140010AAFFE8BFFFFD17DEBA5D002ABFFA2D16AAAA55517D",
INIT_30 => X"020BAFFD17DE10005568B55FF80154BAA280020BA082E82155AA802AAAAFF803",
INIT_31 => X"43FF55085140145F78028BFF08003DF45FFD57FE00FFAABFF45AA803FFEF5500",
INIT_32 => X"842AB55A28015545A284000BA5D53421455504021555D556AB555D5568A00AA8",
INIT_33 => X"2AA800AAAAD142155F7D57DF45FF8002010557FEAAAAF7AABFEAA5D5568ABAA2",
INIT_34 => X"000000000000000000000015555A2FBD75FFA2842ABFF5555575FF55557FEAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000023FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B83008481800E0000C26426040000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"00080D4912E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"000048048002400048150000000002504230C899109032100020160880223000",
INIT_05 => X"040B2A229100410041088011100022201200012840440000B01088C0005C2400",
INIT_06 => X"287E4003225021C5021880C02000A40249048363A5992808110010090908022A",
INIT_07 => X"4044222987020C80152D8910210A0400252B74200045C86810000C5B0503286A",
INIT_08 => X"26509804400501400242C0B0B83B0134702000000000191FA162841324832069",
INIT_09 => X"3002000220001240820F8B2A08000040409018401001200159D80D64AA004041",
INIT_0A => X"020808852000420718C00101B0070310200008B60A23A51B2802467327200801",
INIT_0B => X"080802500C08832582810240812040912094068010050402214850444091019B",
INIT_0C => X"761B011986695014A96E1A8119865A5018C5A0A00012004104020808B0003000",
INIT_0D => X"AE1A811986695014A96E1B0119865A5018C5AF0062C38A4DB680A0D8241501D5",
INIT_0E => X"802CAB184E8F4101621B1BAC845542056A289A1BB2078A922DA2A8B180A2600A",
INIT_0F => X"392000224ACDE215883078681B5C05AA429189B60AC43CEC7F0272C3841DB528",
INIT_10 => X"51BCA1C90006C0C2958502861120C003104289A668B8CAB270106338317A3D94",
INIT_11 => X"A64090B89E015AAA880E48382EB8804B020A06020C67061BC785938085134CD5",
INIT_12 => X"C6284B2D20410AB4503089C00A8280819A5539D503336D61056ABA006282806C",
INIT_13 => X"060040142020015001004A00080042004000E8089C9003066E03513E41470126",
INIT_14 => X"4536708201C000908020349320008000A1000C09A9348498B000000000000080",
INIT_15 => X"32A0C32A0C32A0832A0C19504195040040000000801010028001400010010CBA",
INIT_16 => X"8104400000904C0C0964200841010954000444D280140050C32A0832A0C32A08",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090246811",
INIT_18 => X"1004010040100401004010040102409024090240902409024090240902409024",
INIT_19 => X"0000000000004010040100401004010040100401004010040100401004010040",
INIT_1A => X"488292A831308E0000000A11100830181621409A14E871104201400284000000",
INIT_1B => X"0000000000000000000000000000000000000000000000020820820820820A05",
INIT_1C => X"0000000402000000000000000000010080000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8C0F00000000",
INIT_1E => X"555FFF784020AAF7D542155F7D1400AAF7FFFDE00F7842AA00002A8000000000",
INIT_1F => X"A800AA007FFDFFFA28428A000000001FF08557DF4555516AA00007BEABEFAAD1",
INIT_20 => X"FBEABEFA2D1400AA5D2AAAA00F7FFEAA10F7D17FFFFAAAEA8ABAFFD17FEBAFFA",
INIT_21 => X"0043FFEFA2FFFDE1008556AB45555568A10A2FFC00AAF78028AAAFF84020AAFF",
INIT_22 => X"FFD1555FF0804000AA000428A10AAAA801EFFFD140010AAD57FF45A2D56AA000",
INIT_23 => X"FA2FBFFF550000020000000021EFAA843DE00F7803FEBAFFFFC2000557FC0155",
INIT_24 => X"00F7FBFDEAA007FEAB45AAAE800AAF78428B45A28428A10087FD7400552EBDFE",
INIT_25 => X"A101C2A80000000000000000000000000000000000000000000028BFF5D04154",
INIT_26 => X"AA381C75EABEFBED1575C7E380000BAF7DB4016DE3DF450AAF7F1FDE38FF8A2D",
INIT_27 => X"AFABAFFDF7AE82F7AA870AA0071F8FFFBE842DA101C0E001EF085F7AF6D55556",
INIT_28 => X"42DAAAE38A02082E3FBEFBC7A2DB400824120ADA38E3F1EFA28F7DF7DFD7A2A4",
INIT_29 => X"DF7AF6DB6D56FA3814003AFFFA2F1F8E381C516DB455D5B68A28A2FFC20AAEB8",
INIT_2A => X"BFFC20285D75C2145F7DF525EF140A050AA1C0028A28AAA4801FFE3DF40010AA",
INIT_2B => X"007FD74284120BFFFFBEF1F8F7D080A02038000A001C7A2803AE38FF843DEBAE",
INIT_2C => X"000002DBEF550412428F7F5FDE920875E8B45BEA0850BAE3802DB6DAA8A28A00",
INIT_2D => X"AAF7D57DEAAF7AABDE10552E8000000000000000000000000000000000000000",
INIT_2E => X"1FF007BE8BFF5D516AABA5D5568BEFF7D157555AA80020BAFFFBC01EFA2FFD74",
INIT_2F => X"FEAAF7FBFDF45AA803FEBAFFFBEAA00F7AE974BA085568BEFF7803FE10552E82",
INIT_30 => X"EAAAAA2FFC00AAAA803FEAAA2AA82000A2FFFDF55A2FBC201008003DEAAA2D57",
INIT_31 => X"0001FFAAFFC0010AAFFE8BFFFFD17DEBA5D002ABFFA2D16AAAA55517DF55557F",
INIT_32 => X"802AAAAFF803DEBAAAFBC20BA555142155F7FFC01EF552E974BA550028ABAA28",
INIT_33 => X"2803FFFFA2AAAAA00007FD74BA08003DFFFFFD16ABFF082E820BA082E82155AA",
INIT_34 => X"00000000000000000000003FFEF5500020BAFFD17DE10005568B55FF80154BAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000200000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702684000000008000008820009280A553231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"421A0A0012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"02004000890200001837830011998C31C09060DC104000102002140900003548",
INIT_05 => X"0402002BC200009841090001200006200800000020480010A4100100001C2000",
INIT_06 => X"287FC003230001D0001806C0060CB0622000037085C820000000100C0C200008",
INIT_07 => X"CE64B663DFA314C803292140890C0601F472D1640051F80C10020C493F033432",
INIT_08 => X"67C081000111814004C20481A92940EA7A3020480000071F846890162E135038",
INIT_09 => X"240048108488024082488BAF08000020800629441004300421800F04F8000001",
INIT_0A => X"A0200E0BF40063FF9DC0010000180018200408B27E234913E900067F04D40C01",
INIT_0B => X"002002801000A04200000000000000000000029D204B7C0382FD0100F3F9F80F",
INIT_0C => X"7E0B348EDAC3900F6EFA0B158EDA93900F6EE230381208008001007A80001100",
INIT_0D => X"CA0B158EDAC3900F6EFA0B348EDA93900F6EE8421392C96B1237E0D8BD9628F9",
INIT_0E => X"412EDD2B47CFF812A383430C669E622DBC31D73F6006A5891533EF9500EAE64B",
INIT_0F => X"BA30E022DAD8C100CA39E8CEBE66C2B083798D341B10DE7E14400392C74CAEAD",
INIT_10 => X"71A9C5DD00B12728D5360234D62A49FAB442994B3238D4E2FB104636652E19B8",
INIT_11 => X"C800DA550C29F36A8A2554E48A6430469392526208C6CC95C33717D885329664",
INIT_12 => X"51B60585A5C28895962502E9F36A828C4999AF580395542D27CDBA0020F0FABA",
INIT_13 => X"0000001E404011F066000A000EE040000000873FB80B8A00EF03F56CC12B416A",
INIT_14 => X"4D667C06CC6816B300403C13E2000000460010400000010CE080801010000080",
INIT_15 => X"72F0C72F0872F0872F0C597863978421040800209010124ACA03414158228430",
INIT_16 => X"00104280A89A4D004000000800001D5E05182493C5BC5AF0872F0C72F0872F08",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000010000",
INIT_18 => X"8020080200802008020080200800000000000000000000000000000000000000",
INIT_19 => X"0000000000000080200802008020080200802008020080200802008020080200",
INIT_1A => X"E02000028DCA05A8A28A2048C1111026C152A2316246000CB054420210100000",
INIT_1B => X"C864321904104104104104104104104104104104104104124924924924924481",
INIT_1C => X"2C964B2592C964B2592C964B2592C964B2592C964B2592C964B2190C86432190",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800FFD64B259",
INIT_1E => X"2AA00002AAAA10FF8002155F7FFC2000080417555FFAA80155F7840000000000",
INIT_1F => X"FE8AAA080000155F7FFFDEAA0000020AAF7D542155F7D1400AAF7FFFDE00F784",
INIT_20 => X"2E801FF08557DF4555516AA00007BEABEFAAD1555FFF7842AB55080000145557",
INIT_21 => X"07FFDFFFA28428A00000028B4555043DFFFFFAE82000FF80020AAA2AAAABFF00",
INIT_22 => X"A284174AAFF8428AAAFF8415545AAFBD7545F7AAA8ABAFFD17FEBAFFAA800AA0",
INIT_23 => X"5F7FFFDEAA08556ABEFA2D1400AA5D2AAAA00F7FFEAA10F7D17FFFFAAAE80000",
INIT_24 => X"10A2FFC00AAF78028AAAFF84020AAFFFBC21550800000105D55400AA082A8215",
INIT_25 => X"145F7840000000000000000000000000000000000000000000002AB45555568A",
INIT_26 => X"50AAF7F1FDE38FF8A2DA101C2AAFA00EB8E0516DE3F5C000014041256DEBA487",
INIT_27 => X"2FB551C0E0516D417FEDA921C000017DEBF5FDE92080E000BAF7DB4016DE3DF4",
INIT_28 => X"0070BAAAAAADBD70820801EF085F7AF6D55556AA381C75EABEFBED1575C7E380",
INIT_29 => X"DF7AE82F7AA870AA0071F8FFFBE842DA101C0E2DB55410A3FFC7F7A087000FF8",
INIT_2A => X"7DF7DFD7A2A480000BE8A17482F78A28A92E3841556DA2FBD7545F7AAAFABAFF",
INIT_2B => X"41554508208208017DF7F5FDE9208556FBC7A2DB400824120ADA38E3F1EFA28F",
INIT_2C => X"000002DB455D5B68A28A2FFC20AAEB842DAAAE38A02082E3FBC217D1C0E05000",
INIT_2D => X"005504001FFAA8015545F7800000000000000000000000000000000000000000",
INIT_2E => X"0BAFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE10552EBDE00AAAE975FFAAD1420",
INIT_2F => X"8BEFF7D157555AA803DF45552E975EF007FFFE005504001FFAAD17DE00082E82",
INIT_30 => X"BFF55FF8017410FF84154BAAAAABFF450000021FF007BE8BFF5D516AABA5D556",
INIT_31 => X"BD5555F7AEBFEBAFFFBEAA00F7AE974BA085568BEFF7803FE10552EBDF45002E",
INIT_32 => X"003DEAAA2D57FEAAF7FBFDF45AA8002000FFAE95400F7AEA8A10A284175FFAAF",
INIT_33 => X"2FFC21EF552A954100851554000004021FFFFD17DE1008517DF55A2FBC201008",
INIT_34 => X"00000000000000000000003DF55557FEAAAAA2FFC00AAAA803FEAAA2AA82000A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00020201926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"00104884880A4400403000004800027102A0E88110D83210642EA809C0203040",
INIT_05 => X"04092A08138041184109C001380000201A008128044E00754010C9C192D82400",
INIT_06 => X"201800012372A1D72A180000204024024954A3670819290951001009092C0222",
INIT_07 => X"4000220B40020C80052C0A12292A040005715540015E006810001C4B01032C7E",
INIT_08 => X"9032881000140140024200808839005C002010800000155F8122851320016400",
INIT_09 => X"2C80080200801280825A988008000040008208401005B3071859006442004054",
INIT_0A => X"200810940400720005C0030192072310200028B6022346080802E001A5600801",
INIT_0B => X"206822F20CA8826AC2A14250A128509528954404144C200425010040000001B0",
INIT_0C => X"A41AA5B7344C10B383081BA4B7341C10B3831034081200000000000430003000",
INIT_0D => X"381BA4B7344C10B383081AA5B7341C10B383110218CB0E54C2EA404A4F03D404",
INIT_0E => X"A008E730A01AB113A5524E6ACA678001CE3E20A5B284ED1132909C72885A2B2C",
INIT_0F => X"6430202021252991C22C99731014AC3CC0C0B8182597A801610218CB0C3548B3",
INIT_10 => X"5194332B018A444AEA2701288A15A151EC5952E44128CA194517354C180A3C06",
INIT_11 => X"D50048A411C158BB0A7910142C771804C8A0ADA2E6A983014780CA28B2A5C882",
INIT_12 => X"F8BE8E3E1E0109472C3EB50158BB02D09852745F80112C428562EE0353635232",
INIT_13 => X"02414032646000826080C20001104240480068001C9B9150A0000297046E4023",
INIT_14 => X"4510008241C80290882400908000A000A1000809A93485D61000000000000080",
INIT_15 => X"00000000040000000000000020000000000000008010102A82014100101118BA",
INIT_16 => X"A10441010090480C096420184321040002844840000000004000000000400000",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094246A10",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"0000000000005094250942509425094250942509425094250942509425094250",
INIT_1A => X"BFBFBFBF7DDF3BAAAAAABEFDDFE7EFBEFFE7CFC3F7EFFF7DF7E24502A8000000",
INIT_1B => X"F5FAFD7EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAFFD",
INIT_1C => X"BF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EB",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800FFDFAFD7E",
INIT_1E => X"80155F7842AB55552E821FFFFD5555EF552ABDFEF007FE8A00AAFBC000000000",
INIT_1F => X"BD55EFAAD1554BA00556AA00AAD16AA10FF8002155F7FFC2000080417555FFAA",
INIT_20 => X"55420AAF7D542155F7D1400AAF7FFFDE00F7842AA00002A821EF5D7BC21FFFFF",
INIT_21 => X"80000155F7FFFDEAA00002AB45082A821EF5D557FF45A2AABFEBA082A975555D",
INIT_22 => X"A2FFE8BEF5D517FF455D554214500043DEBAAAFFEAB55080000145557FE8AAA0",
INIT_23 => X"0552EBFEAAAAD1401FF08557DF4555516AA00007BEABEFAAD1555FFF7842AABA",
INIT_24 => X"FFFFAE82000FF80020AAA2AAAABFF002E80000AAAABDF555D2E955EFA28428A1",
INIT_25 => X"A28AAF5C0000000000000000000000000000000000000000000028B4555043DF",
INIT_26 => X"000014041256DEBA487145F78428B6D4120851FFEBD5525C74124B8FC71C71EF",
INIT_27 => X"871C74975C01FFEBF5D25EFA2D555482085F6FA28AAD16FA00EB8E0516DE3F5C",
INIT_28 => X"0BFE921C2E9557D415B400BAF7DB4016DE3DF450AAF7F1FDE38FF8A2DA101C2A",
INIT_29 => X"0E0516D417FEDA921C000017DEBF5FDE92080E2AB7D1C24851FF495F7FF55A2A",
INIT_2A => X"ED1575C7E38028A82B6F1E8BFF495F78F7D49554214508003FEAABEFFEFB551C",
INIT_2B => X"5D20905C7AA842DA00492EBFEAABED1401EF085F7AF6D55556AA381C75EABEFB",
INIT_2C => X"000002DB55410A3FFC7F7A087000FF80070BAAAAAADBD7082087000AAA4BFF7D",
INIT_2D => X"4508042AB455D517DEBAA2D54000000000000000000000000000000000000000",
INIT_2E => X"E00AAAE975FFAAD1420005504001FFAA8015545F78028BFF0004175EFA2D5421",
INIT_2F => X"DEAAF7AABDE10552E975450051401EFA2D5421EFAAD557410007BFDEAAA2D57D",
INIT_30 => X"175FF087BFFF45AA843FE005D2A955FF087BC20BAFFFBC01EFA2FFD74AAF7D57",
INIT_31 => X"03FEBAFFFBFDF45552E975EF007FFFE005504001FFAAD17DE00082EA8BFF5504",
INIT_32 => X"516AABA5D5568BEFF7D157555AA8028A00FFD16ABFF087BEABEF005542155000",
INIT_33 => X"00017410AA803DFEF550402155A2843FE00082ABFEAAFFD5421FF007BE8BFF5D",
INIT_34 => X"00000000000000000000003DF45002EBFF55FF8017410FF84154BAAAAABFF450",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000033FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"0002074F200904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000480488024000403000000000001002A0E881108032100002000800203040",
INIT_05 => X"04092A081000411841080001000000201000012800400010001081C000402000",
INIT_06 => X"80500001221021C1021800002000240249048361001128081100100909000222",
INIT_07 => X"4000220050020480152D0A142D0A8400043B45400040006810000C5901033D78",
INIT_08 => X"0010880000100140024280808829029C002000000000053FA142051324902030",
INIT_09 => X"2000000000000200820888800800004000800840100020011858006442004040",
INIT_0A => X"200800840400400005C0010190070310200008B202236D080802400001600801",
INIT_0B => X"000000100C088020028102408120409120940404104C20002101004000000110",
INIT_0C => X"5210040000B0E0A0000210040000E0E0A0000190081200000000000000003000",
INIT_0D => X"0210008000B0E0A0000210008000E0E0A0000B02740421A0E5D1A02400205080",
INIT_0E => X"40110080A4006110510C14D18178E01200860008920106460D4501CB00011130",
INIT_0F => X"411420220080220C0093C38923240ABBC00905C33C6000400F02740412C0715C",
INIT_10 => X"8000120800658992F3C700C3018120000041DB011CC000090012565306500002",
INIT_11 => X"E240240A8340000200067EAA8CB65809240C09024A4AE0CA0000480083968239",
INIT_12 => X"7DB0D0200900422ACA4B28000002002B46867DBC002A830280000800F7B7A0B1",
INIT_13 => X"020040126060008020000200000042004005800004801150A00341244000845C",
INIT_14 => X"4500008240800000802000908000800001000009A92481041000000000000080",
INIT_15 => X"000040000000000000040000000000000000000080101000000141001001088A",
INIT_16 => X"810440000090480C096420084101040000044040000000004000040000000000",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090246810",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"0000000000004090240902409024090240902409024090240902409024090240",
INIT_1A => X"EFBBBBAABCDABF9E79E7BEF9CB91FE1EF7D3AEB9F3E6FF7DF650400280000000",
INIT_1B => X"FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7FC",
INIT_1C => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8FF000FE7F3F",
INIT_1E => X"E8A00AAFBE8BEFA2D568ABA00003DF555555574AAAAAEAAB45082E8000000000",
INIT_1F => X"02AABA555155400557BC2010557BEAB55552E821FFFFD5555EF552ABDFEF007F",
INIT_20 => X"002AA10FF8002155F7FFC2000080417555FFAA80155F78428AAA007FE8A10080",
INIT_21 => X"AD1554BA00556AA00AAD140145AA8028ABA002EBFFFF082EBDEBAA2D1420105D",
INIT_22 => X"A2AEA8A10080428A10FFAEBFFEF5D0428B45A2FFC21EF5D7BC21FFFFFBD55EFA",
INIT_23 => X"5F7FBC0010FFAA820AAF7D542155F7D1400AAF7FFFDE00F7842AA00002A80155",
INIT_24 => X"EF5D557FF45A2AABFEBA082A975555D55400BA005568A000000175FFF7D15554",
INIT_25 => X"B6D00248000000000000000000000000000000000000000000002AB45082A821",
INIT_26 => X"25C74124B8FC71C71EFA28AAF5E8BFFB6D56DA82000E38F6D4155504AAA2AEAA",
INIT_27 => X"28ABA147FEDA10080E2AAAA555552400417FC20005D75E8B6D4120851FFEBD55",
INIT_28 => X"4BAEAAB6DB4202849042FA00EB8E0516DE3F5C000014041256DEBA487145F784",
INIT_29 => X"75C01FFEBF5D25EFA2D555482085F6FA28AAD147155BE8028A82002EB8FC7002",
INIT_2A => X"F8A2DA101C2A80145B6AEA8A10080E2DA00F7A0BDFD7550428B55A2F1C71C749",
INIT_2B => X"0004175FFE3D15757DE3F5C0038FFAA800BAF7DB4016DE3DF450AAF7F1FDE38F",
INIT_2C => X"000002AB7D1C24851FF495F7FF55A2A0BFE921C2E9557D415B400AA00556DA00",
INIT_2D => X"EF0051400AAA2AAAABFF08000000000000000000000000000000000000000000",
INIT_2E => X"BFF0004175EFA2D54214508042AB455D517DEBAA2D568BEFFFD57FE10002AAAB",
INIT_2F => X"01FFAA8015545F78028AAA557FFFE00082EAAAAA5D5142000007BC20105D5568",
INIT_30 => X"28A00082EAAB45000028ABAFFFBC20AA08043DE00AAAE975FFAAD14200055040",
INIT_31 => X"02AB55AAD1575450051401EFA2D5421EFAAD557410007BFDEAAA2D557555FF80",
INIT_32 => X"FFD74AAF7D57DEAAF7AABDE10552E82155FFAAA8A10002ABFE00F7803FF555D0",
INIT_33 => X"87BC20AA00517DE000804175EFAAD1555EFA2D1420BAFFAE820BAFFFBC01EFA2",
INIT_34 => X"000000000000000000000028BFF5504175FF087BFFF45AA843FE005D2A955FF0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000100000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"000440009282000001100000000000100220C8811080321000000228002A3000",
INIT_05 => X"04092A0010004300418800510000A6201000012A64400000145080C000422000",
INIT_06 => X"00100001220001C00018821020402402080003772019200001001009090002AA",
INIT_07 => X"4000220000021840010C8912250A0400042044400040006810000C4901032B18",
INIT_08 => X"0022810000058140024280A0A8190004002030C00000016F8122041320000000",
INIT_09 => X"20000000000002C0820888008800000000800840100020011850004402004040",
INIT_0A => X"00080094000062000180010180060210200008B2022304080800400003E00801",
INIT_0B => X"0000000008008020020000000000000100800000000000002500004000000130",
INIT_0C => X"0010108000000000000010108000000000000230001200000000000420003000",
INIT_0D => X"0010140000000000000010140000000000000100000040000000000000000000",
INIT_0E => X"0000000000000100008040000000000000000000020000090000000000000000",
INIT_0F => X"0030002000406000000000068409014000000000000000000100000040000000",
INIT_10 => X"0000000800000201000800000000000000400048000000000010000440000000",
INIT_11 => X"00A0000000000002000000441108800000000002008008000000000080201000",
INIT_12 => X"0242038B82800000000000000002000001000000000000000000080000001844",
INIT_13 => X"000000100000000005C04A000000400000000000000001062000000400000000",
INIT_14 => X"4500008200800000800000100000800001000001A12480001000000000000080",
INIT_15 => X"000000000000000000040000200002000000000080101000004140001001088A",
INIT_16 => X"0004400000904808094020080000000000044040000000004000040000400004",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000046000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000400280000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000000000",
INIT_1E => X"AAB45082EBFE000004020AA552E80000F7FBC214555003DE10A2FBC000000000",
INIT_1F => X"BE8A10F7802AA0055003FE10007BE8BEFA2D568ABA00003DF555555574AAAAAE",
INIT_20 => X"AEAAB55552E821FFFFD5555EF552ABDFEF007FE8A00AAFBFDEBA555568BEFA2F",
INIT_21 => X"55155400557BC2010557BFFFEFA2FFC20005D2A955EFF78428BEFAAD17DF55AA",
INIT_22 => X"5D2AA8B45AAD57FF55A2FBC21FFA28415400FF8028AAA007FE8A1008002AABA5",
INIT_23 => X"A002E9740055516AA10FF8002155F7FFC2000080417555FFAA80155F7843DF45",
INIT_24 => X"BA002EBFFFF082EBDEBAA2D1420105D003FFFF08514200055002AA00AA802AAB",
INIT_25 => X"E28B6FFC0000000000000000000000000000000000000000000000145AA8028A",
INIT_26 => X"8F6D4155504AAA2AEAAB6D0024B8E381C0A00092412A87010E3F5C0145410E3D",
INIT_27 => X"F8EAA495F68BFFA2F1EFA38E38428A005D0038E28147FE8BFFB6D56DA82000E3",
INIT_28 => X"428BEFB6DB7DF45AAAEA8B6D4120851FFEBD5525C74124B8FC71C71EFA28AAF5",
INIT_29 => X"7FEDA10080E2AAAA555552400417FC20005D75F8FFFBEF5C0000492A955FFF78",
INIT_2A => X"BA487145F7843FF7D4120A8B6DAAD17FF55B6F5C21EFAA8E10400E38E28ABA14",
INIT_2B => X"41002FA38A2842AA82142095428415F6FA00EB8E0516DE3F5C000014041256DE",
INIT_2C => X"0000007155BE8028A82002EB8FC70024BAEAAB6DB4202849043FFC7005F45010",
INIT_2D => X"00A2D542155002ABDEBAF7FBC000000000000000000000000000000000000000",
INIT_2E => X"BEFFFD57FE10002AAABEF0051400AAA2AAAABFF08002AAAA5D2A82000082E954",
INIT_2F => X"AB455D517DEBAA2D56AABA087BEABEFAAD57DEAAA2802AA105D002AABA5D7BE8",
INIT_30 => X"42010082A955EFFF8428BFFFFFBFDF55A2AEA8BFF0004175EFA2D54214508042",
INIT_31 => X"A82000AAAAA8AAA557FFFE00082EAAAAA5D5142000007BC20105D556ABFFF7D1",
INIT_32 => X"D1420005504001FFAA8015545F7803FFEF08002ABEFA2D57DF45F7D1401FFA2A",
INIT_33 => X"8043FF55087BD740000043DEAAA2842AA005D00154AA007BFDE00AAAE975FFAA",
INIT_34 => X"000000000000000000000017555FF8028A00082EAAB45000028ABAFFFBC20AA0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000300000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"0202115002BB10080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"2FE962000017102918900948514522CE09200C0D590569398ADBF8CC1E50E480",
INIT_05 => X"5E6023002834854AE41C1E8782F508F2A15B71D412E0AFD9C2990DA56FF0B55A",
INIT_06 => X"B9B9E55402000340003200220A86012D0000000480D0400001555960540180A0",
INIT_07 => X"40D890101DBD400901442800817C2901F400868554DE240000A80090CE82A803",
INIT_08 => X"0122004000005665510320C9C90510025A8A00000A0A048F550A440E0001380C",
INIT_09 => X"2060410280081116C8204D016CB2CB290008008279580411289000000118A905",
INIT_0A => X"00008176802203180025699200140001A15000017F0051D0F837324E002A8A56",
INIT_0B => X"4485D000000124002400000000000001004010A8812831605DA0000A054052E4",
INIT_0C => X"B5320018CAC99BA0A3B9320018CAAAADA0C343F1AC1B01040A00202489551455",
INIT_0D => X"59320018CAC99BA0ACB9320018CAAAADA0CC421CA003B694B68018FAAA708E2C",
INIT_0E => X"B2449A3FF2FA04E5E09B128834ADB1443A1891E4A928C29020E6A8524CE7A3EE",
INIT_0F => X"2375B801324301AB0067622E5E5404B2A5A40B1E6644AF0F021EA003AC24352A",
INIT_10 => X"0A8C241815FEB6A9158863F638FB60ED838E890B703C6260D8E3A21275714C90",
INIT_11 => X"15F11133D171727A2550EE2F1BA0064F70DBDB1C74424E91E1C194C71D1216F5",
INIT_12 => X"432A2B2D001F803471A9A960E57245FDF9D364DBD9435A6D45C9E81BED555E4C",
INIT_13 => X"C00006B0800000038814B72AB01508150013F162119014204373517700ACCC59",
INIT_14 => X"300208092B940192D1000000000000A8A5AA80018120E00066000000000012CA",
INIT_15 => X"1000110001100011000108000880008000520228080108039501200848002912",
INIT_16 => X"081500008A422150884081AC9000010003561180063DB4F61100011000110001",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000012000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"BCBF0F2C688A8D3CF3CF0A7A898D21B4C9838D3030EF5168A360400000000000",
INIT_1B => X"E9F47A7D345345345345345345345345345345345345345145145145145147A5",
INIT_1C => X"3E9F4FA3D1E8F47A3D1E8F47A3D1E9F4FA7D3E9F4FA7D3E9F4FA7D1E9F47A7D1",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800001F4FA7D",
INIT_1E => X"3DE10A2FBC21FFFFFBFDF45A2D56AB45FFFFD54BAFF80001FF002A8000000000",
INIT_1F => X"FFFE005D7BC0010002E954AA087FFFE000004020AA552E80000F7FBC21455500",
INIT_20 => X"FFE8BEFA2D568ABA00003DF555555574AAAAAEAAB45082E974BA5D7BFDF55A2F",
INIT_21 => X"7802AA0055003FE10007BC0000082A97400550017410FFD1555550000020BAAA",
INIT_22 => X"AAFBD74105504021FF5D2EAAABAFFFBD55FF002ABDEBA555568BEFA2FBE8A10F",
INIT_23 => X"0007FC00AA087FEAB55552E821FFFFD5555EF552ABDFEF007FE8A00AAFBD55EF",
INIT_24 => X"005D2A955EFF78428BEFAAD17DF55AAAE820AA5D517DF45AAFFFFEAAFFAABFE1",
INIT_25 => X"1FF08248000000000000000000000000000000000000000000003FFEFA2FFC20",
INIT_26 => X"7010E3F5C0145410E3DE28B6FFC21C7E3F1F8F55AADB6FB6DFFFBD54AAE38E02",
INIT_27 => X"92482497BFDF45AAFFF8E385D7BC5000002E904BA1C7FF8E381C0A00092412A8",
INIT_28 => X"B555450804070BABEF5E8BFFB6D56DA82000E38F6D4155504AAA2AEAAB6D0024",
INIT_29 => X"5F68BFFA2F1EFA38E38428A005D0038E28147FC2010142E90428490015400FFD",
INIT_2A => X"C71EFA28AAF5D25D7B6F1D54384904021FF5D2AADAAAFFF1D55FF002EB8EAA49",
INIT_2B => X"A2F1FDEAAEBAABDE001471C20921475E8B6D4120851FFEBD5525C74124B8FC71",
INIT_2C => X"0000038FFFBEF5C0000492A955FFF78428BEFB6DB7DF45AAAE820925D5B7DF45",
INIT_2D => X"EFF7FFD54AAAAAA801EF00000000000000000000000000000000000000000000",
INIT_2E => X"AAA5D2A82000082E95400A2D542155002ABDEBAF7FBC2145AAD568B45AAFBFFF",
INIT_2F => X"00AAA2AAAABFF080000000087BFDF55A2FFE8AAA557FD7410082A800AA557BEA",
INIT_30 => X"800BA080417400F7FBD75450800174AAFFD168BEFFFD57FE10002AAABEF00514",
INIT_31 => X"1575EF082EAAABA087BEABEFAAD57DEAAA2802AA105D002AABA5D7BC20005D2E",
INIT_32 => X"D54214508042AB455D517DEBAA2D540155F7D1554AA0800001EF5D2ABDEBAF7D",
INIT_33 => X"2AE82010557FFDF55A2D57FEAAAAAEBFE10555140000555568BFF0004175EFA2",
INIT_34 => X"00000000000000000000002ABFFF7D142010082A955EFFF8428BFFFFFBFDF55A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000100000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"5295B6957FCBE0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"6DE90201BF90102103AF158E805428249851BFB2C106592088DBF8400A5055C2",
INIT_05 => X"3824BD7F80148D9E07100A8201ED01C1A19B68F40A807ED9C18114956FF081DB",
INIT_06 => X"6A8F033DD800000000050716BE9F57F8AC000807DFD9B00000CF20E5E1818B1B",
INIT_07 => X"86481240FE05A109228E2C0891D772A6F40045B8CF30E085DD2ED57D4EED08CA",
INIT_08 => X"DF23800005981C0338190549C904182B6113870022000488C08B46268A001508",
INIT_09 => X"823DF78CDB6CA60E0E28EFFE2061872F80C1684A80C8604085F0074D3B72637F",
INIT_0A => X"BD2FAD7FE653C3BA1FF33E0E001E000B3A5DAADAFDDA5DA79350CFB8013E7437",
INIT_0B => X"C5C3D00018006C681700000000000000020012E9E10A31EB5FF9296A67F5B4FF",
INIT_0C => X"542A6FEEB2533EA160782A6FEEB2333EA16031F2BD47BDA2CA5D8164FCCFE833",
INIT_0D => X"F82A6FEEB2533EA160782A6FEEB2333EA160391BEFF2C32FB695F919110D5ECE",
INIT_0E => X"5A86840354D1706FFFA3EF6E24B6D18C0D06638A207CFDE1F7DDAD76D5282400",
INIT_0F => X"4D77FAAB77CE3AF3EE78F58DB737E6E43E59AFE4A59B57679D19EFF2C7573FAD",
INIT_10 => X"72CA52606DFED6CA55334C04C04FF7D7A0ABD6DAAAB96529382B74E4E1FE4ACA",
INIT_11 => X"AA1A184045D5D7A870D2F5A5D7522D1281017F056E9C9C3FC95949C157ADB555",
INIT_12 => X"A58949D5B5C85F97871876F7D7E859FDEB974F486905001FDF5FA0D719F9956E",
INIT_13 => X"70021EE341036BF368128419FB5560158015177F916A039EF41FDB34A91F432E",
INIT_14 => X"1D0A7CC9AE7A08BFF0001D35682AC0CE8FCCC200A59BDD2FFE3F3EC7C7DEF206",
INIT_15 => X"BCF4FBCF4FBCF4FBCF4FBE7A7DE7A7800617112E46F05D02DD814102F800633F",
INIT_16 => X"00179C16DECF67F08BC02F9086000D9E8A3F06ABD73DBCF4FBCF4FBCF4FBCF4F",
INIT_17 => X"000000000000000000000000000000000000000000000000000000000005F080",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"930D0D1B9000303AEBAE88BE013DB9880A5D25C0408006114F981800C0000000",
INIT_1B => X"351A8D069A6BAE9A69A6BAE9A6BAE9A69A6BAE9A6BAE9A69A69A69A69A69A918",
INIT_1C => X"A351A8D46A351A8D46A351A8D46A341A0D068341A0D068341A0D068351A8D068",
INIT_1D => X"00000000000000000000000000000000000003FFFFFFFFFFFFFF8000011A8D46",
INIT_1E => X"001FF002A821FFFFFFFFFFFFFFBFDFEFAAD142010007BEAB55FFAA8000000000",
INIT_1F => X"A975EFA2D140145007BC21FF5D2A821FFFFFBFDF45A2D56AB45FFFFD54BAFF80",
INIT_20 => X"7BFFE000004020AA552E80000F7FBC214555003DE10A2FBEAB45A28000010082",
INIT_21 => X"D7BC0010002E954AA087FD7400082E954AA0800154AA0855575FFAAD57FE005D",
INIT_22 => X"F7D16AB45FFFFEABEF007BD74005555555EFF7AE974BA5D7BFDF55A2FFFFE005",
INIT_23 => X"5555568B45552EA8BEFA2D568ABA00003DF555555574AAAAAEAAB45082EBFFFF",
INIT_24 => X"00550017410FFD1555550000020BAAAFFC0145AA84154BA082E801FFAAFBC015",
INIT_25 => X"B7DEBA480000000000000000000000000000000000000000000000000082A974",
INIT_26 => X"FB6DFFFBD54AAE38E021FF0824851FFFFFFFFFEFF7F1FAFD7A2D5400001C7BED",
INIT_27 => X"EFB45AA8E070281C20925FFBEDB451451C7BC01EF4124821C7E3F1F8F55AADB6",
INIT_28 => X"5505EFBEDB7AE385D7FF8E381C0A00092412A87010E3F5C0145410E3DE28B6FF",
INIT_29 => X"7BFDF45AAFFF8E385D7BC5000002E904BA1C7FD54280024924AA1404174AA005",
INIT_2A => X"2AEAAB6D0024BFFD7FFDB6AB7DFFF5EDBC71C7BD54005D5B575EFEBAE9248249",
INIT_2B => X"1C20801FFB6F5C0145555B68B7D4124A8BFFB6D56DA82000E38F6D4155504AAA",
INIT_2C => X"0000002010142E90428490015400FFDB555450804070BABEF5C516DAA8A12492",
INIT_2D => X"45AAD5400005D7BFFFEFAA800000000000000000000000000000000000000000",
INIT_2E => X"145AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF0000155FFF7FBFDFEFFFD568B",
INIT_2F => X"2155002ABDEBAF7FBFDF55A2AA974AA5D04001EFFFFFD5545557BC21FF080002",
INIT_30 => X"000AA5500174AA0855421FFFFFBEAAAA5D7BEAAAA5D2A82000082E95400A2D54",
INIT_31 => X"BD75FFAAAA80000087BFDF55A2FFE8AAA557FD7410082A800AA557BD74BA0004",
INIT_32 => X"2AAABEF0051400AAA2AAAABFF08003FF55F7FFEABFFF7D57FF455D7FD54105D7",
INIT_33 => X"FD1555FFA2AA800105504001EFFFD140145557BE8BEF000028BEFFFD57FE1000",
INIT_34 => X"0000000000000000000000020005D2E800BA080417400F7FBD75450800174AAF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000033FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"080BA868803F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"42016B0C401F58495C900A4859552A611D9A640F5903B2388004004C08A06008",
INIT_05 => X"16226B107811422A641C08038040007060E0032801E0202000991B708280B501",
INIT_06 => X"B3B8E0FC86142B4142B0000000011114D305824024090A1A143F182000000000",
INIT_07 => X"802102401015610A02C4005000EA019D002482043FCF1C8090C02800C0120886",
INIT_08 => X"20D40A5004003260F9810541494D403D9B98810A0002C601000054B94A006880",
INIT_09 => X"6070000504102805C820C8016C30C250080C0182183804012A0A102200110180",
INIT_0A => X"E000108010230445A800FD865421432121804021C20452880C2D100000022E0C",
INIT_0B => X"C2060014250B9080008306C18360C1B0609C05013065CC042004040808084001",
INIT_0C => X"8582081483ACC15F9C3982081483CCC15F9CBA45505640000A402019003F140F",
INIT_0D => X"F982081483ACC15F9F3982081483CCC15F9FB1962FCB69E08AAAEAEBCDDF7C72",
INIT_0E => X"E3F8E7F5E3AC3620805298B15A3FEBF1CFFF7670ACC3811A28AB57523CDFEBFB",
INIT_0F => X"DC4041D4CF03138DD865103EFEEAC9002BF05800D875E63CC9962FCB52CAA02F",
INIT_10 => X"8DB7BFE25208E8F46A228BF8A757F1B72A8A800B7546DB9F1CA320037F01BD67",
INIT_11 => X"9509EAAE7FD3B749471C48F8A45981CCFAFDBF9464006FD037AEFAE5150016EA",
INIT_12 => X"8802A3AF8E8FB0440CE78773B709641256EC844B8AF92FD7CEDC24A9E181A8A2",
INIT_13 => X"C284601C2864000080113307E4800297D086E00036D2440E0880AAD62BEFF577",
INIT_14 => X"A88DCC2211E44174112840880000060D7030C30B885200D274004008080003C1",
INIT_15 => X"0308003080030800308001840018400400602A01880980037109700C04C44C92",
INIT_16 => X"8340000020301805002D008CD943626111C0D95C20C2030A0030800308003080",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B0680834",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"00000000000041B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1",
INIT_1A => X"60B22A145DF60B8208209679D701DC2E784601F95163897DF160000000000000",
INIT_1B => X"944A2512AAA8A28A28A2AAAAAA8A28A28A2AAAAAA8A28A28A28A28A28A28A244",
INIT_1C => X"8944A25128944A25128944A25128944A25128944A25128944A25128954AA552A",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8000004A2512",
INIT_1E => X"EAB55FFAA821FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E820BA55000000000000",
INIT_1F => X"16AB55A2D542000A2D5400BA0800021FFFFFFFFFFFFFFBFDFEFAAD142010007B",
INIT_20 => X"80021FFFFFBFDF45A2D56AB45FFFFD54BAFF80001FF002A821FFFFFFFFFEFF7D",
INIT_21 => X"2D140145007BC21FF5D2AAABFFF7D168B45AAD57DFFFFFFFC0010F7842AA10F7",
INIT_22 => X"000002010552E95410AAFBD75FF5D7FEAB5500516AB45A28000010082A975EFA",
INIT_23 => X"5A284155FF5D517FE000004020AA552E80000F7FBC214555003DE10A2FBEAA00",
INIT_24 => X"AA0800154AA0855575FFAAD57FE005D7BD74000804174AA5D00020BA55554214",
INIT_25 => X"0AA490A00000000000000000000000000000000000000000000017400082E954",
INIT_26 => X"AFD7A2D5400001C7BEDB7DEBA4871FFFFFFFFFFFFFFFFDFEFF7FFD74AA552A82",
INIT_27 => X"821FFF7F1F8FC7EBD568B7DB6DF47000AADF400AA080A051FFFFFFFFFEFF7F1F",
INIT_28 => X"1C2000F78A2DA38E38A021C7E3F1F8F55AADB6FB6DFFFBD54AAE38E021FF0824",
INIT_29 => X"8E070281C20925FFBEDB451451C7BC01EF4124ADBC7E3D56AB7DB6DF78FD7EBF",
INIT_2A => X"10E3DE28B6FFE8A101C0E05010412495428AAF1D25EF497FEAB7D145B6FB45AA",
INIT_2B => X"5D0A000BA555F47145BE8A105EF555178E381C0A00092412A87010E3F5C01454",
INIT_2C => X"00000154280024924AA1404174AA0055505EFBEDB7AE385D7FD7438140012482",
INIT_2D => X"EFFFFBD54BA5D2A820AA082A8000000000000000000000000000000000000000",
INIT_2E => X"5FFF7FBFDFEFFFD568B45AAD5400005D7BFFFEFAA80155FFFFFFFFFFFF7FBFDF",
INIT_2F => X"54AAAAAA801EF0000021EFF7D16AB55A2D56ABEFF7FBD5410AAFBC00AA002A95",
INIT_30 => X"68BFFF7FFEAB45AAD140010F7AABFEBAAAAA82145AAD568B45AAFBFFFEFF7FFD",
INIT_31 => X"BE8BFF557BFDF55A2AA974AA5D04001EFFFFFD5545557BC21FF08003FF55AAD1",
INIT_32 => X"2E95400A2D542155002ABDEBAF7FBE8A00552E954100000154AAA2D1421FF007",
INIT_33 => X"D7BD74BA5D0002010552E820AA5D7BD7545F7AA801EF55516AAAA5D2A8200008",
INIT_34 => X"0000000000000000000000174BA0004000AA5500174AA0855421FFFFFBEAAAA5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000100000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000010228001000000000000000000024001620280000000000354200004008",
INIT_04 => X"00016200001310090090004840004152C7208802590000388000004C08006000",
INIT_05 => X"1621008008100002641C0803804000702000000000E02000009900000000B100",
INIT_06 => X"0210200C00000000000000000000000080000000000000000003182000000000",
INIT_07 => X"C00D267001B880080700285020020AC98820022802400480405008901100A001",
INIT_08 => X"000000000000106009872048400C4000010D000008000204150A00815A010084",
INIT_09 => X"0000000000000004C80000002C30C200000000021808005800000000000E0E00",
INIT_0A => X"0000000000000000080025860000000080A00020602040800000000000022A04",
INIT_0B => X"C002000000000000000000000000000000000000000000000000000084000760",
INIT_0C => X"385598035D0008A003B05598035D0008A0034078104B41A41000000000031400",
INIT_0D => X"505598035D0008A000B05598035D0008A0004263C0343EDD414004042228DC0D",
INIT_0E => X"0401180DE053A98F6ECC739D8140040231068187C39F5A4F985C008902041124",
INIT_0F => X"227848D4303807FC8CC5508AEAED1BFBD406451B02000E033263C0343CB74050",
INIT_10 => X"00000018A700FCF980CC300318A2420851546B2400000040D8549B5800000010",
INIT_11 => X"40E40511802208D6B30C48F8A8A452210402120A936B0000000004C2A8D64800",
INIT_12 => X"0006362A2B6424287B08286208D6B1427ED430B41402D025082359700181C211",
INIT_13 => X"40000000000000000010030060009C000018440021011821B35254E99AF9E941",
INIT_14 => X"002000044000000000000000000002F0001F00002024B20002000000000002C0",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000040",
INIT_16 => X"00000000000000000000008C8000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"441189B9045D82A69A69803F47E18E0218CC0140400200441920000000000000",
INIT_1B => X"4C261309861861861A69861861861861A69861861861861861861861861861A1",
INIT_1C => X"84C26130984C26130984C26130984C26130984C26130984C261349A4C2613098",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000261309",
INIT_1E => X"820BA55003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A800105D2E8000000000",
INIT_1F => X"FFDFEFF7FFD54BA5D2EA8BFFFF84021FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E",
INIT_20 => X"AE821FFFFFFFFFFFFFFBFDFEFAAD142010007BEAB55FFAABDFFFFFFFFFFFFFFF",
INIT_21 => X"2D542000A2D5400BA08003DFFFFFFFFFFFFF7FBE8B55A2D540010007BEAABAA2",
INIT_22 => X"FFFFFDFEFA2D56AB45AAFBD74AAFFD5420100804021FFFFFFFFFEFF7D16AB55A",
INIT_23 => X"AFF802ABFFFFAE821FFFFFBFDF45A2D56AB45FFFFD54BAFF80001FF002ABDFFF",
INIT_24 => X"45AAD57DFFFFFFFC0010F7842AA10F780155FFF7FBE8B45AAD568BFFF7FBD74B",
INIT_25 => X"000412A8000000000000000000000000000000000000000000002ABFFF7D168B",
INIT_26 => X"DFEFF7FFD74AA552A820AA490A38FFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2A80",
INIT_27 => X"BAFFFFFFFFFFFFF7FBFDFD7EBF1D24AA5D2AADBD7E384071FFFFFFFFFFFFFFFF",
INIT_28 => X"140000007FEFA92A2AA851FFFFFFFFFEFF7F1FAFD7A2D5400001C7BEDB7DEBA4",
INIT_29 => X"F1F8FC7EBD568B7DB6DF47000AADF400AA080A3FFFFFFFBFDFC7E3F5EAB45AAD",
INIT_2A => X"38E021FF0824BDFEFE3F1F8FD7AAD16DB7DBEFBD74AAE3DF400000004021FFF7",
INIT_2B => X"B6DB6FBD7E3F5D04AAFF8A2DBD7E3A0821C7E3F1F8F55AADB6FB6DFFFBD54AAE",
INIT_2C => X"000002DBC7E3D56AB7DB6DF78FD7EBF1C2000F78A2DA38E38A125C7E3F1EAB55",
INIT_2D => X"FFF7FBD54BA552A80010002A8000000000000000000000000000000000000000",
INIT_2E => X"5FFFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA082AA8BFFFFFFFFFFFFFFFFFF",
INIT_2F => X"00005D7BFFFEFAA8028BFFFFFFFDFEFF7FFFFF55A2D5400AA552ABDF55A28015",
INIT_30 => X"FDF55AAD16AB55AAD140010007BFFE10AAAA955FFF7FBFDFEFFFD568B45AAD54",
INIT_31 => X"BC20100800021EFF7D16AB55A2D56ABEFF7FBD5410AAFBC00AA002ABDFEFF7FB",
INIT_32 => X"FBFFFEFF7FFD54AAAAAA801EF00003FFEFA2D56AB45A2D57DFFFFFFFD54AAA2F",
INIT_33 => X"AAA82155AAD568B55FFFFFDF55A2D1400AAF7AABFF45AA8002145AAD568B45AA",
INIT_34 => X"00000000000000000000003FF55AAD168BFFF7FFEAB45AAD140010F7AABFEBAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000200000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"0001E6000053300B00D0005800000000000000407B0004BB830004DC3D01E000",
INIT_05 => X"FEE0000008720043EC3C3D0F87FA19F7E0201C409BE1F10623BB000A100CF300",
INIT_06 => X"06102FFC8E0007C00078008000171175A200096404D9404003FFDBE4744200AA",
INIT_07 => X"482491301000010001DC00000000000000004203FE4005800000008030002000",
INIT_08 => X"20E2008000027FEFF946058180010429000001080AAA010F8000000000000000",
INIT_09 => X"400000120000913FD80000003DF7DE0080010047FBF8000000000800C5408000",
INIT_0A => X"0080000010000400080FFDBE000000400000010000010050600220461003EAFE",
INIT_0B => X"C00600000000801020000000000000010240001721214E000004000000080000",
INIT_0C => X"08020000200000000F30020000200000000F3008001E00000000001803FF14FF",
INIT_0D => X"F0020000200000000F30020000200000000F3040200000020000000026A70C00",
INIT_0E => X"000019B140000800800000020000000030B86000400080000200000000004A58",
INIT_0F => X"AC08000000508001030A0A4001000000000002183E61E6000040200001000000",
INIT_10 => X"0000A56000090100000000001F86C00010080000000000525801000000000014",
INIT_11 => X"0000001716800000803102020000000002BC360020000000000292C010000000",
INIT_12 => X"DF70C08040100000706707600000801000000000000057450000100106060000",
INIT_13 => X"C011001C81080001101F977FE00800000000000040040040002000080506049C",
INIT_14 => X"0000000000000000020020029000000000000000020000000000000000000ADF",
INIT_15 => X"0000000000000000000000000000000000000000000002000200000000000000",
INIT_16 => X"0801810100000000000093ED8000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000401008080",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"930424038000343CF3CF349600704000201120A983400E0104D2040020000000",
INIT_1B => X"190C86432CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB0C30C30C30C30C818",
INIT_1C => X"2190C86432190C86432190C86432190C86432190C86432190C86432190C86432",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8000010C8643",
INIT_1E => X"800105D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8201008040000000000",
INIT_1F => X"FFFFFFFFFBD54BA552A8001000003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A",
INIT_20 => X"2E821FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E820BA5500001FFFFFFFFFFFFFF",
INIT_21 => X"7FFD54BA5D2EA8BFFFF843FFFFFFFFFFFFFFFFFFFFEFF7FFD74BA552E801FF00",
INIT_22 => X"FFFFFFFFFFFFBFDFEFFFD542000082EAAB55AAAABDFFFFFFFFFFFFFFFFFDFEFF",
INIT_23 => X"0087BE8B55F784021FFFFFFFFFFFFFFBFDFEFAAD142010007BEAB55FFAA801FF",
INIT_24 => X"FFF7FBE8B55A2D540010007BEAABAA2AE975FFFFFFFFFFFF7FBFDF55AAD14000",
INIT_25 => X"00014000000000000000000000000000000000000000000000003DFFFFFFFFFF",
INIT_26 => X"FFFFFFFBD54AA5D2A80000412ABFFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A82",
INIT_27 => X"021FFFFFFFFFFFFFFFFFFEFF7FBD74BA5D2A800281C0038FFFFFFFFFFFFFFFFF",
INIT_28 => X"FD54BA5D2A801C7142E871FFFFFFFFFFFFFFFFDFEFF7FFD74AA552A820AA490A",
INIT_29 => X"FFFFFFFF7FBFDFD7EBF1D24AA5D2AADBD7E38438FFFFFFFFFFFFFFFBFDFEFFFF",
INIT_2A => X"C7BEDB7DEBA4871FFFFFFFFFEFF7FBF8FD7E3D140010142AAFB7DBEAEBAFFFFF",
INIT_2B => X"E3F1FAF45A2D142010087FEDB55F78A051FFFFFFFFFEFF7F1FAFD7A2D5400001",
INIT_2C => X"000003FFFFFFFBFDFC7E3F5EAB45AAD140000007FEFA92A2AA925FFFFFFFDFEF",
INIT_2D => X"FFFFFFD74AA552A820005D040000000000000000000000000000000000000000",
INIT_2E => X"BFFFFFFFFFFFFFFFFFFFFF7FBD54BA552A80010002ABFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"54BA5D2A820AA082A821FFFFFFFFFFFFFFBFDFEFF7FFD74AA5D2A800BA550428",
INIT_30 => X"FFFEFF7FBFFFFFF7FBD74BA552A80145552E955FFFFFFFFFFFF7FBFDFEFFFFBD",
INIT_31 => X"ABFFFFFFAEA8BFFFFFFFDFEFF7FFFFF55A2D5400AA552ABDF55A2802ABFFFFFF",
INIT_32 => X"D568B45AAD5400005D7BFFFEFAA80175FFFFFBFDFEFF7FFEAB45AAD1420105D2",
INIT_33 => X"AAA821EFF7FBFDFFFAAD168B55A2D542010007BFDF55F7AE955FFF7FBFDFEFFF",
INIT_34 => X"00000000000000000000003DFEFF7FBFDF55AAD16AB55AAD140010007BFFE10A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"1094EC681244819000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"0001E6000053300F01D4587800446194F49020107F0012BBC00202DC3823EA82",
INIT_05 => X"FFF201B228704123FC3C381F87C03DFFF012412A9FE1E01013BF09404050F300",
INIT_06 => X"96F43FFF002004020044041084CB01AD000003761702401000FFDFE050000080",
INIT_07 => X"043C802A821D41412001A0040950AB60014114C3FE4187A009A663A680100B30",
INIT_08 => X"2C01004000047EFFF811A46968004060629A0002208A00000068113205A12034",
INIT_09 => X"0A812D8D5B742D3FF84056383FF7DE0880042107BFF9C45B85101C49A37F4000",
INIT_0A => X"0822189000480406310FFDFE00040009814C089202225412115414601DE3EBFE",
INIT_0B => X"C0281280080180B2948004400220011100841200D001000624000100C002804A",
INIT_0C => X"60694101816002D41A4068C101815004D8158809C86065941840B1014FFF56FF",
INIT_0D => X"0068C101816002D41A40694101815004D815810D42E04A08A80098C024500253",
INIT_0E => X"12682960828F05C96A001B029010134160C8125B0B271802242880A04482418A",
INIT_0F => X"100920C54E8EA256ECF078BA081C10080E05C0B06AA8B12CFD0D42E0441A3000",
INIT_10 => X"4F30A8801406D00290006280320100010362A8A20826A88660D86B202049F115",
INIT_11 => X"2011819E290048A2118EC8140C08064802C0081B0D64040936443306C5514410",
INIT_12 => X"C40A0300600C0A80509F418008804581BA0038005A706680012280506A801060",
INIT_13 => X"C000120080002341881F3FFFF80DCC158092C044600466208CC5091011C322A4",
INIT_14 => X"398C6021569249C4B3007127080806FF917FC30010107688862A28C54518DBFF",
INIT_15 => X"228D9228D9228D9228D99146C9146C84006309044081A001B188300E20806520",
INIT_16 => X"8004000000E07008010003EF80022A51904595123203040D9228D9228D9228D9",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010044800",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"0000000000004010040100401004010040100401004010040100401004010040",
INIT_1A => X"FFBFBFFF7CFE7F9E79E7FFEDDFEFFFBEFFE7DF83F7EFFFFDF7E0000000000000",
INIT_1B => X"FDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FBFDFEFF7FB",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800003FFFFFF",
INIT_1E => X"8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8001000040000000000",
INIT_1F => X"FFFFFFFFFFD74AA552E80010552EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A",
INIT_20 => X"2ABDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A800105D2EBFFFFFFFFFFFFFFFF",
INIT_21 => X"FFBD54BA552A800100000001FFFFFFFFFFFFFFFFFFFFFFFBD54BA5D2E8201000",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF7FBD74BA5D2E800BA5D00001FFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A552A800BA5D2E821FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E820BA5500001FF",
INIT_24 => X"FFFFFFFFFEFF7FFD74BA552E801FF002E975FFFFFFFFFFFFFFFFFFEFF7FBD74A",
INIT_25 => X"00008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA552A8200014003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E80",
INIT_27 => X"BDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2E800005D2ABFFFFFFFFFFFFFFFFFF",
INIT_28 => X"BD54BA552E82028002AB8FFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2A80000412A",
INIT_29 => X"FFFFFFFFFFFFFFEFF7FBD74BA5D2A800281C00001FFFFFFFFFFFFFFFFFFFFF7F",
INIT_2A => X"52A820AA490A071FFFFFFFFFFFFFFFFFFEFF7FBD74AA5D2E800AA5500021FFFF",
INIT_2B => X"FFFFFDFEFF7FFD54BA5D2E80082492E871FFFFFFFFFFFFFFFFDFEFF7FFD74AA5",
INIT_2C => X"0000038FFFFFFFFFFFFFFFBFDFEFFFFFD54BA5D2A801C7142E955FFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8000008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005D043FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"54BA552A80010002ABDFFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2E800005D2EBF",
INIT_30 => X"FFFFFFFFFFDFEFF7FBD74AA552E820BA002AA8BFFFFFFFFFFFFFFFFFFFFF7FBD",
INIT_31 => X"E800BA5D04021FFFFFFFFFFFFFFBFDFEFF7FFD74AA5D2A800BA5504021FFFFFF",
INIT_32 => X"FBFDFEFFFFBD54BA5D2A820AA082A955FFFFFFFFFFFFFFBFDFEFFFFFD54BA552",
INIT_33 => X"52E975FFFFFFFFFEFF7FBFDFFFFFFBD74AA5D2E80000082A955FFFFFFFFFFFF7",
INIT_34 => X"00000000000000000000002ABFFFFFFFFFEFF7FBFFFFFF7FBD74BA552A801455",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"8632CA211E4491D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"24B000808800040439245B221373581F97B0A8D1040F92000F42000047A00E58",
INIT_05 => X"011B2BBA308F023810004700083E220811E9BF2844021B1004045E4249500449",
INIT_06 => X"80A51003AA0200C020088E16A85235722940A817251101010100040D6D0702A2",
INIT_07 => X"5C9ECAB0D247B013B405EAD525FAE48FC2060B880081A26DCD4047EFF9EF0189",
INIT_08 => X"2D0141C0055280100751096B6A40D6F86723E510AA2004803D3275EB2024E814",
INIT_09 => X"04804818CD280100207246A8020000AC0283002004051507A5411C0DA0005048",
INIT_0A => X"2C6898B2950AA65635B00041C23020131A80CFDFF3FE509A907C556828201102",
INIT_0B => X"050F60E220A06880D2A14050A028501428054278142151262CA50343854E506A",
INIT_0C => X"612B3482C0C0078E1F412B1582C090078E1F840A2B0114020104022460002200",
INIT_0D => X"012B1582C0C0078E1F412B3482C090078E1F891C239F8908003099C1ACF06273",
INIT_0E => X"1BA859F213AFC14AA380430060181BA1B0FD16770236A4091621C08055C2C0DB",
INIT_0F => X"B08AA600CA88B143AB11880C280600101F09C030AB28B03C111C239F87082804",
INIT_10 => X"4B61BD8068B92400D0004E30368910E8822A984B0025B0DE6089462660095337",
INIT_11 => X"001AC2173B00E162563454C40804055412D4481128C4CC012A66F30455309600",
INIT_12 => X"50840180A00E1C81900C4190E160589C48082C006A9057CA4385809520F07830",
INIT_13 => X"004416B105036B4180C000800C8C00460848952220592745AC11A544B1BF0068",
INIT_14 => X"512C6A8C4F0008AA800470370000A0004D0000002126F30C902A29C54539C020",
INIT_15 => X"2A81C2A81C2A81C2A81C9540E1540E001400006100003202D040050220103D2A",
INIT_16 => X"22365034A8EA754008004C0214202C50013456520CA09281C2A81C2A81C2A81C",
INIT_17 => X"104411044110441104411044110441104411044110441104411044110445E220",
INIT_18 => X"0401004010040100401004010040100401004411044110441104411044110441",
INIT_19 => X"0003FFFFFFFF9004010040100401004010040100401004010040100401004010",
INIT_1A => X"FFBFAFBEFDFFBBBEFBEFBEFBDFD1FE3EFBD7ADF9B3EFDF7DF7D0512289000000",
INIT_1B => X"FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79EFFC",
INIT_1C => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000FE7F3F",
INIT_1E => X"8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2A8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8201008043FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74AA552E80010552EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E8000055",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD54AA5D2A82000552ABFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2A800005D2EBDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A800105D2EBFFFF",
INIT_24 => X"FFFFFFFFFFFFFFBD54BA5D2E82010002AA8BFFFFFFFFFFFFFFFFFFFFFFFFD54A",
INIT_25 => X"0100004000000000000000000000000000000000000000000000001FFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001008043FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74AA552E800105D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A820001400",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD54AA5D2E800005D2ABFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A80000412AB8FFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A82010552EBDFFFFF",
INIT_2B => X"FFFFFFFFFFFFBD54BA552E80038492EB8FFFFFFFFFFFFFFFFFFFFFFFFBD54AA5",
INIT_2C => X"00000001FFFFFFFFFFFFFFFFFFFFF7FBD54BA552E82028002AA8BFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201000040000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74AA552A820005D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001000043F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD54AA552E8001055003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"A820105D2ABDFFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2E800005D2EBDFFFFFFF",
INIT_32 => X"FFFFFFFF7FBD54BA552A80010002AA8BFFFFFFFFFFFFFFFFFFFFF7FBD54BA5D2",
INIT_33 => X"02AAABFFFFFFFFFFFFFFFFFFEFF7FBD74BA552E800AA082EA8BFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000000021FFFFFFFFFFFFFFFFDFEFF7FBD74AA552E820BA0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"5886C0201A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"0005EE040057700F40D08078500000D9218020407F0000BB8018A2FC380BEAC2",
INIT_05 => X"FFE0419028700023FCBC385F87C0BFFFE0124002FFE1E0C517FF09111212F300",
INIT_06 => X"16D03FFC96102081020000020489019C430480241202080810FFDFE000000000",
INIT_07 => X"0001160A003475C8100123400E20E1F40F439647FF4807E189A477EF81DF0AF1",
INIT_08 => X"801008000007FEFFFB110140695812CC4188D58A0AAA10803448D0844FB71000",
INIT_09 => X"4201258112D4487FF8001010FFF7DE4000000003BFF8C25818080020017F0F94",
INIT_0A => X"0C024000004A9400000FFDFF50010103134CAFDF03BA18000F39900037C3EBFD",
INIT_0B => X"C02812F00429DC92C40002000100008000105400C00400100000A01800080100",
INIT_0C => X"A1CAF13F214001521001CBF03F21100152100801C17E61841950B1C10FFF57FF",
INIT_0D => X"01CBF03F214001521001CAF13F2110015210088528E00E02C8200A430A424202",
INIT_0E => X"02C86040902AC60BACDF0E02D02001C1C044006D0C94FB94320880603C420B80",
INIT_0F => X"00010AF5052419D196441902801430182800A018D9CA8000648528E00D124802",
INIT_10 => X"4D101808458A5602E000892029110445C19960A00026880C006739000009B003",
INIT_11 => X"1009408021144CB042F880100C0601844068880CE72000013600600332C14000",
INIT_12 => X"F80E02120018390320F050144CB241D0B9023402085020825132C8CB5B404030",
INIT_13 => X"C200400020224000405F7FFFE0008E17C0D240406519400500840A9524EE38A1",
INIT_14 => X"AC810033149249C433200180082A06FF907FC308181204800600000000001BFF",
INIT_15 => X"010C1010C1010C1010C10086080860840063090442A18001B188300C48907120",
INIT_16 => X"0100000000000004002403EFC10302219A41C1443243050C1010C1010C1010C1",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200010",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000080200802008020080200802008020080200802008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000000000",
INIT_1E => X"8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8001000043FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2A8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA552A8200000043FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A552A8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8201008043FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74AA552E8000055003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2A8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E800000800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA552A8001008043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52A8200014003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8200008043FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74AA552E820101C003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E800105D043FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000043F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2A8001008043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"A8200008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001000043FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74AA552A820005D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552",
INIT_33 => X"5003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA552E8200055043FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA552E800105",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"0000745C200801000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"0001E6000053300F00D0007810042140C00000407F0000BB800000DC3801EA00",
INIT_05 => X"FFE0000008700003FC3C380F87C019FFE01240009BE1E00003BF00000000F300",
INIT_06 => X"06103FFC000000000000000004890088010080001202000000FFDFE000000000",
INIT_07 => X"0009B24B043980021000810284204A8001401643FE4007E5501AA00000DC8C30",
INIT_08 => X"0000000000007EFFFB11A56940581280031D61420000B080102040BC5B006120",
INIT_09 => X"020125811254083FF80000003FF7DE0000000003BFF8005800000000017F0000",
INIT_0A => X"0000000000000000000FFDFF4000000AA0354000019C40000128000011C3EBFC",
INIT_0B => X"C000104000000010440000000000000000001000C00000000000000240058000",
INIT_0C => X"4012500021B00880108012500021E00880104809C1666594584031010FFF56FF",
INIT_0D => X"0012500021B00880108012500021E0088010492064206100E81084200048C080",
INIT_0E => X"0410004C840041A0D8005410903804100144800803419043064900C002050184",
INIT_0F => X"020902F60002260D65B361BAA1041018140F02C0000809408D20642053027004",
INIT_10 => X"00020818B06D9802F00030C02060110002C9E8010C00010480B35A0300400041",
INIT_11 => X"20042108603100061516EE800C060228204300166B4060080008240593D00218",
INIT_12 => X"7C02000040206602C10B48110006143B62023C00142800B04400095DFF902030",
INIT_13 => X"C000000000000000001F17FFE000DC1180C7804400044029208301040214AE4C",
INIT_14 => X"008000010012414433000100080806FD107FC300000000000600000000001BFF",
INIT_15 => X"000C1000C1000C1000C100060800608400630104408180012188300C00814080",
INIT_16 => X"0000000000000000000003EF80020201904181003003000C1000C1000C1000C1",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"F30C2416857732AEBAEBFFA55EDCF9822659AE7BE742E6441990000000000000",
INIT_1B => X"3C1E0F07BEFBEFBEF9E79E79E79E79E7BEFBEFBEFBEFBEFBE7BE7BE7BE7BEC98",
INIT_1C => X"83C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F078",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8000001E0F07",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008040000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8001000043FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2A8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008040000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2A8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008040000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8000008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000043FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8000008043FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A800100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00004000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"4909E6093253306F82D0007C80000000080E01007F8020BBC00040DC3801EA00",
INIT_05 => X"FFE0000008704503FE3C380F87C019FFF01241009BE1E00203BF80800000F392",
INIT_06 => X"06103FFF9E2086C2086E006604C9019D03108B741202605040FFDFE070400880",
INIT_07 => X"4024057000000100000000000000000001401643FE4007C00000000000CC0830",
INIT_08 => X"0801404000007EFFFF40010000401408000045000000A0801000408000000000",
INIT_09 => X"4A7DF795965C6D3FFC0020003FF7DF01880C618FBFFDD75E00100040437F0000",
INIT_0A => X"0000000000009400000FFDFFC006020000000000019804000028000191C3EBFF",
INIT_0B => X"C02812E0182000F2C48304418220C11160845004D04820000000000000000000",
INIT_0C => X"0002400001000800000002400001000800000801C0786184185031810FFF56FF",
INIT_0D => X"0002400001000800000002400001000800000000202000000800000000080080",
INIT_0E => X"0000000404000000880000001000000001000000000090000008000000040000",
INIT_0F => X"000100C600800001040000040009100000000200200000400000202000020000",
INIT_10 => X"0002000000081001000000000040010000082000000001000001080000000040",
INIT_11 => X"0080000040010000001080001008000000010000210000000008000010400000",
INIT_12 => X"0000030280000000010000010000001020000000000000100400000108000040",
INIT_13 => X"E0120012C1400080291F17FFF0018C11808200400000400000C2000000042000",
INIT_14 => X"00800001001243443B000100880806FD107FC301800000000600000000001BFF",
INIT_15 => X"000C1000C1000C1000C10006080060840077330C4889CC292588300C00804000",
INIT_16 => X"82068C0200000008014023EF80020201904189003003000C1000C1000C1000C1",
INIT_17 => X"110441104411044110441104411044110441104411044110441104451044C820",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FFFFFFFFFFFFC110441104411044110441104411044110441104411044110441",
INIT_1A => X"200A625D144BC2B4D34D7F61432D518B45265EF8278C2015DA080800002FFFFF",
INIT_1B => X"88C4623124924924924924924924924904104104104104104124904124904281",
INIT_1C => X"58AC562B158AC562B158AC562B158AC562B158AC562B158AC56231188C462311",
INIT_1D => X"00000000000000000000000000000000000003FFFFFFFFFFFFFF800002C562B1",
INIT_1E => X"8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"0003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"94A7B2B1450000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"6FEBEF5FEC737AFBC6F85FDEB220109E1FEFFFE3FBA7FDFB9BD301DC3FF5F0D2",
INIT_05 => X"FEEDBFDC387F987FEF7C3FAF87FF59F7F5FB7FF59BE1FF980BBBB7FE6D21F3DB",
INIT_06 => X"57902FFDEE9D7DC9D7DF2B263893479DDFAFDFE15213FEFEBFFFFBE1F1D3A333",
INIT_07 => X"10992310605CE10301DE0C1831CB7DF60A244B9BFEE00589DDBCEFEDC1DFA089",
INIT_08 => X"001D8EA111DA7FEFF90F21C8C84D9C0D858FC7020828C18FD18346BBF0000180",
INIT_09 => X"F37DF7B9DF7DCB3FDE89ECC07DF7DF5F985C6BCFFBFA28F99E7EB07F47FFEFAA",
INIT_0A => X"7DCFE1D4077B4D0026FFFFBE7D67D7F3BB79CFFB83BF14EC1E7D5980580BFAFF",
INIT_0B => X"C7D7D51D6F5FDCB935D7AFEBD7F5EBFBF7FEBD66DBFCA3F87501AE7B08060730",
INIT_0C => X"01F45EC0010007E01001F45EC0010007E010084BCD7FF1B61B5C33813FFFFCFF",
INIT_0D => X"01F45EC0010007E01001F45EC0010007E01001BD8020500008001F0100405202",
INIT_0E => X"1EC00040B02007EC09A0E00010001DC0004600400F781429C0080000770001A0",
INIT_0F => X"404B3BFD0402346235408402C08010003C064000E408010081BD802060020000",
INIT_10 => X"0E401A08FE0012040000FC002001360403E434588007200D00F88C84C081C203",
INIT_11 => X"001F01002156040675809145400007B00040091F1190982038406807C868B100",
INIT_12 => X"008320C0403C34000088601604067D00212000007C400082D81009FC08281D00",
INIT_13 => X"F7BFFED3FBFF6A84383F177FF005FFBFF5FA1040076065F730FC08043A903A80",
INIT_14 => X"F589807B7096CD4CF73AC1FC98884FFF19FFC71FEFED7B251E35768E8ED6BFDF",
INIT_15 => X"8C0D78C0D78C0D78C0D7A606BC606B8C56F7730ECCDBDF152199F51EDDCDEBCF",
INIT_16 => X"DFE7DD87FEFF7FF796FFFFFDFFD7E681B867D3683A03A40F78C0D78C0D78C0D7",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFEFDFD",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"FFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEB",
INIT_1A => X"57AA9ABAD8ACBF0E38E3A89F9E923C2CD990A7D0D2A377F86EDB5C88646FFFFF",
INIT_1B => X"4C261309861861861861861861861861861861861861861861A69A6986186EBC",
INIT_1C => X"84C26130984C26130984C26130984C26130984C26130984C26130984C2613098",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000261309",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"1085B0B041000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"6FAB975B6470BAF386C87A9CB00000001FEF9F23E3A7BDE79B5101D23FB5C0C2",
INIT_05 => X"F8EDBFD4347F18778E723F2E47FE59C7F5FB7F759B91FB880BA3B6FE2921CBDB",
INIT_06 => X"47000FFC128D5CE8D5CC210638A046889CAB57E8421786B6ACFFE3E181932377",
INIT_07 => X"000000042000000288020C18300320620A80231BFE200181092CE7ED80DFC001",
INIT_08 => X"000C562551D87E8FF90041101042110180004102800008801183468180000141",
INIT_09 => X"137FF7A0FF75813F1C85244071EFBF17D85C738BE3FA08F9DE36B05B07FEEF22",
INIT_0A => X"768EA0C406630D00226FFE3E2D62D6E21259CFDB039E806C02451880400BE0FC",
INIT_0B => X"CC57550D63564D1D2556ADAB56D5AB6AD7EAB962CBD8A3A83101F47E08040510",
INIT_0C => X"01E44A40010007600005E44A4001000760000843C561E5C55C42B9011FFF48FF",
INIT_0D => X"05E44A40010007600005E44A40010007600004BD8020100008001F0100001302",
INIT_0E => X"1EC00000382006EC0820A00010001DC0000208400D781020C008000077000020",
INIT_0F => X"40431BC50402146235400400408010003C064000C400018080BD802020020000",
INIT_10 => X"0E400204FE0010040000FC0000003E0403A424108007200102E888808081C200",
INIT_11 => X"001F0100005E040475808101400007B00000015D111010203840081748482100",
INIT_12 => X"00012040403C34000080201E04047D00202000007C400000F81001FC08080500",
INIT_13 => X"E5ADA4C25ADE72041A3F147FF0018DBBB5FA10400360649310FC08003A903A80",
INIT_14 => X"054880693016DD4C755AC16C1A884FFE18FFD757E7ED7A211E81C09818109E1F",
INIT_15 => X"440C3440C3440C3440C3C2061A2061AD46FF730E5CCBCD55219AB55F0DEFABC7",
INIT_16 => X"5EC71385FC2512E3565BBBF1BAD6F281BC63F1683803C00E3440C3440C3440C3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BDE75ED",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"FFFFFFFFFFFFAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB",
INIT_1A => X"200E5E48710A4200000028150200903950C086D0E28028104A471688747FFFFF",
INIT_1B => X"0080402000000000000000000000000000000000000000020800000000000780",
INIT_1C => X"5028140A05028140A05028140A05028140A05028140A05028140201008040201",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8000028140A0",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"8C2100804900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"02000100440408002408008002221000204116A280000F000001400000100010",
INIT_05 => X"0004D44400004D4400000000000000000000005C0000000A0000002C20600000",
INIT_06 => X"4100000120040A0040A00B0090006202940100004000A2020400200888800911",
INIT_07 => X"5002489020420110800244891211440804000810002000081040000000200000",
INIT_08 => X"080542C004CA00000050080202008401842004108AAAA00008912240A1248804",
INIT_09 => X"0000000C0000E400002040500000009202C1002040004400022200020400B062",
INIT_0A => X"58C460540329810002D002000400407020800000004000640800088008280001",
INIT_0B => X"0140000401028008330000800040002002480102010082981500062108020430",
INIT_0C => X"00040A40000000A00000040A40000000A0000040060084104110828030000800",
INIT_0D => X"00040A40000000A00000040A40000000A0000000800010000000000000005000",
INIT_0E => X"00000000A00000040020A000000000000006000000080020C000000000000120",
INIT_0F => X"4040152000000020000004004080000000000000240000000000800020000000",
INIT_10 => X"0000120002000004000000000001220000040410800000090000808080800002",
INIT_11 => X"0000000001420000200001014000000000000900101010200000480008082100",
INIT_12 => X"0001204000000000000820020000200000200000000000028800002000080500",
INIT_13 => X"00933050080C0001900020000000408010000000022000D61028000008000000",
INIT_14 => X"400082D022040000400800081022C0000080000206CB0821082B694D4D294000",
INIT_15 => X"050160501605016050160280B0280B0012000843066021001400040024440245",
INIT_16 => X"0861CD33548542A10209D4100E4040A00002002C004001036050160501605016",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008021081084",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"0000000000000020080200802008020080200802008020080200802008020080",
INIT_1A => X"06A0A0F108816B1861863BED822140048D2E5818732C5589A40A0C22E1000000",
INIT_1B => X"80C0603020820820820820820820820820820820820820820820820820820035",
INIT_1C => X"582C160B0582C160B0582C160B0582C160B0582C160B0582C16030180C060301",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800002C160B0",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0803B2814D0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"26E1E905CC574828C4F85FC600000016004F77E2F887CDB80BC340DC07D1F000",
INIT_05 => X"FE1DFE4C080F884FE33C078F803F19F011E93ED49BE01F1A03B8972E6D20F049",
INIT_06 => X"57902000DE142D4142D5030010134395D70589415002DA4A17FFF800F0C38111",
INIT_07 => X"00092300601CE00101DE040811D919F402244293FEE00400CCB46BA4C164A088",
INIT_08 => X"08148A4000887FE0000F20C8C80D080D818FC2000000418FD08142BAD0000884",
INIT_09 => X"E204D2154D28AA3FC60888D03C10415A80402847F8002458926A002E457FA0AA",
INIT_0A => X"5587A1540231410006DFFF80540541619968C76980E914E4163D4980100BFA02",
INIT_0B => X"07C7C0140D0B50A8218102C0816040B1225C1506512C83E85500AC3A08040630",
INIT_0C => X"00141EC0000000A01000141EC0000000A01008480D3EB4A24A0C910037FFFC00",
INIT_0D => X"00141EC0000000A01000141EC0000000A0100100800050000000000000405200",
INIT_0E => X"00000040B000010401A0E000000000000046000002080429C0000000000001A0",
INIT_0F => X"40483B590000202000008402C080000000000000240801000100800060000000",
INIT_10 => X"00001A08020002040000000020013600004414588000000D00108484C0800003",
INIT_11 => X"000000002156000220001145400000000040090210909820000068008828B100",
INIT_12 => X"008320C00000000000086016000220000120000000000082D800082000281D00",
INIT_13 => X"32936E43A92F2880B01F37001004B29450580000066021F6303C000408000000",
INIT_14 => X"B481806A62840800C22800B8900042FF0180000ABFEF89250815568A8AD6ABC0",
INIT_15 => X"8D0068D0068D0068D006A68034680300021410028450530014014002D445624D",
INIT_16 => X"89418D13FE7F3FFD8BADB7FC4F4164A00806522C0A40A50268D0068D0068D006",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C4B12C9894",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"FFFFFFFFFFFFC0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0",
INIT_1A => X"FFBF3F5E7CFC7DFFFFFFD7FADDCFFFBEFFCF1F879DFFFFFDFFEA0C00602FFFFF",
INIT_1B => X"DFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBAEBAEBAEBAEBAFFFD",
INIT_1C => X"FDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800003EFF7FB",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"F7AEBEBFFDFFBFBEFBEFFFFFDFF3FC3EFFF7FDFBF76FF7FDFFD0000000000000",
INIT_1B => X"FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79EEBD",
INIT_1C => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000FE7F3F",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"1084B030000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"6DA986092050306382C05A1C900000001FAE89016387B2A38B5000D03FA1C0C2",
INIT_05 => X"F8F92B90307F41338E303F0E07FE19C7F1FB7F289B81FB8003A396D20940C3DB",
INIT_06 => X"06000FFC020004C0004C000628800488080003600213001000FFC3E101030222",
INIT_07 => X"000000000000000220000810200220620E00030BFE000181092CE7ED80DF8001",
INIT_08 => X"0000000001107E8FF90001000040100000004102200000801102448100000100",
INIT_09 => X"027DF780DF74013F1C00240071E79F05888C618BA3F800599C101049037E4F40",
INIT_0A => X"240A808004420400202FFC3E002202021259CFDB039E0008024510000023E0FC",
INIT_0B => X"C407500020004C10060204010200810040801060C04821202001A05A00040100",
INIT_0C => X"01E04000010007400001E0400001000740000803C0616184184031010FFF40FF",
INIT_0D => X"01E04000010007400001E04000010007400000BD0020000008001F0100000202",
INIT_0E => X"1EC00000102006E80800000010001DC0000000400D7010000008000077000000",
INIT_0F => X"000308C50402144235400000000010003C064000C000010080BD002000020000",
INIT_10 => X"0E400000FC0010000000FC000000140403A020000007200000E808000001C200",
INIT_11 => X"001F01000014040455808000000007B00000001D010000003840000740400000",
INIT_12 => X"00000000403C34000080001404045D00200000007C400000501001DC08000000",
INIT_13 => X"E004048240426200081F147FF0018C1380DA10400140640100D4080032903A80",
INIT_14 => X"050800A91012494C31004124080886FE187FC301B124F2001600000000001A1F",
INIT_15 => X"000C1000C1000C1000C18006080060840477330C4889CC012188310E08812982",
INIT_16 => X"02061004A820104809402BE1900222019861D1403803800C1000C1000C1000C1",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100446020",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"FFFFFFFFFFFF8100401004010040100401004010040100401004010040100401",
INIT_1A => X"00000000000000000000000000000000000000000000000000001000802FFFFF",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000000000",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"ED39BA795990D275FB4A6E96ACC4731DEA4598B0AFB54867F6EE4618C3749807",
INIT_01 => X"58A0047D8607944AC7DA180001ECA2544042106208408208C20022E9173734B3",
INIT_02 => X"9F775E7CB273E6CCA7DAAF00001000000478020113C9C38E09FB7CCCDD9F203E",
INIT_03 => X"88280C4C7B4CB04443163C91110C58F24A31000B8028A810A3D0F8B169A01006",
INIT_04 => X"00160090920C04800904848262220277E05152B280780D407428E723C01E1400",
INIT_05 => X"0006D46207801E400183C0707800E6000E008057641E00473C40680D32330C00",
INIT_06 => X"C165000225E2C11E2C12A0D0144AC27206582C166504816162002000B0FC21D5",
INIT_07 => X"5E6D233B964E7CD99DFB870E1DDDD889C5FBDC440129A0604442180238203F70",
INIT_08 => X"AD23C17544C581000657A0E8E83D86F0E4A7B2D88AAAFD7FE0E1833AC5920CFC",
INIT_09 => X"6D82082E2081B6C0027ADA398000008A504318404005B70663212C04A080B036",
INIT_0A => X"414568729139FA5610C00001A2502440888420247041E87681008CE9AFC80001",
INIT_0B => X"22B826E250B12346F1244812240912048941621804A150CA1CA45C254D4AF4AA",
INIT_0C => X"F80FA97FE0F0009E0FC40FA97FE0F0009E0FC048211E9C11C31F82E4A0008900",
INIT_0D => X"040FAB3FE0F0009E0FC40FAB3FE0F0009E0FCC42EFDFBF0AE03080E2AEB2E0F1",
INIT_0E => X"013879BA878FE807F65FBF12E0380231F0BD9E3FC08FEBD6F661C0E008C3CB5F",
INIT_0F => X"B248831ACBFC8BBDCAB779BC699F20180309A0F83BE2B87C7C42EFDFBF187806",
INIT_10 => X"4131B59003FFEC07F00003F01FB90BE9F01FC8B38C2098DAE007F323A0C83136",
INIT_11 => X"3080E29F1B2BE9F8A27E6E915C0E004C72BEC800FE7464290626D7003F994718",
INIT_12 => X"FC0C2352A0024B83F07F198BE9F8A0FFDA2A3C0202B8776A2FA7F023F7D06570",
INIT_13 => X"1448126105810941C5C068000CD4004C0905E52630BB1AE49C2BA7F98D6F846D",
INIT_14 => X"6074EA560F0416A24844B01302A26100C4801844069B0C88881A28C141118000",
INIT_15 => X"A781E2781EA781E2781C33C0613C0E21020800239450116ED443C041B47E9665",
INIT_16 => X"241140A056954AB0C280D0002020187007122C3E04E03383E2781EA781E2781E",
INIT_17 => X"20481204812048120481204812048120481204812048120481204812058112C1",
INIT_18 => X"0481204812048120481204812048120481204812048120481204812048120481",
INIT_19 => X"0000000000001204812048120481204812048120481204812048120481204812",
INIT_1A => X"C4109CAF9C4C83B8E38E2AE9C136AD8E9B562CF042E6281CF13043A85D400000",
INIT_1B => X"F0F87C3E08208208208208208208208208208208208208208208208208208220",
INIT_1C => X"1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F87C3E1",
INIT_1D => X"000000000000000000000000000000000000C3007FFFFFFFFFFFA00000F87C3E",
INIT_1E => X"4214555517DEAA5D7BFFEAAF7803FEBAF7FFD74BAAAAABDEBAF7AE8000000000",
INIT_1F => X"1555FF55517FE000055421FF00557DF45A2D5401EFF7D142145A2AE800BA0851",
INIT_20 => X"5555555A2AABFFFF5D516AA00A28028A00AAAEBFE00A2FBD75FFFF8400155085",
INIT_21 => X"5517FF45A2AEBDEBAAAAAA8BFFF7D140010FF84174BA552EBDFFF0004020005D",
INIT_22 => X"5504000BA5D2E97545A28028B4508554014508043FEBA082ABFE10AAAEA8ABA5",
INIT_23 => X"FA2AABFE00FFFFD74AA085540000002E801FF557FD75FF0051401FF5D0015410",
INIT_24 => X"EFF7FFC20BAF7D1575450800020BA08517FF45F7FBFFF45A2FFFDE00002E801F",
INIT_25 => X"A38BF8FC000000000000000000000000000000000000000000002ABEFAA80001",
INIT_26 => X"7155BC2A87092AAFA9257F1C5BC00AA5D7FF8EAA57803AEBAF7F5D74AAA2A03A",
INIT_27 => X"BFBC7EB8005B55A85B555EF095F50578085BE8FC7A3F00516DA2D5451D7EBDB4",
INIT_28 => X"0975FFAAA1521FF492BF8F40B6AAB84AF555168A00EA8000150A801C01C7142E",
INIT_29 => X"2EBAE28168ABAA2D43D568BC5400168E90E2F412BEAE3D542A004380124921D2",
INIT_2A => X"2FA3AA28EA8168A954100071D2E90A855C7A00A38F6DE05B40480557A95A3A1C",
INIT_2B => X"16D1EAE925EA0BFEBF4AA09217F490568417085147B50A80095178157FEFA074",
INIT_2C => X"000002D57AAA8402A8743DBD202DA95568A95E800A8F57F6DA971F8F7FFFA42D",
INIT_2D => X"AAFFD1564BA2282BFA02A2C28000000000000000000000000000000000000000",
INIT_2E => X"5EFA87F57555AAFBD7555FFAE95408A8FDC31AD017D34ABA5D7BEAAAAD786BCE",
INIT_2F => X"C2087383F79A5046A37B55F38415555797D63BFF007F8B2B2D97D483AFA7BD9F",
INIT_30 => X"42000D382964A92B401E71D7581C33172EC0A0300A6AEA8FAF0451CA001D4845",
INIT_31 => X"C8365A2FD5E04AA5780A8AAAD7AC3CA02003BEBBA7D7463CC508D07577BAFBD5",
INIT_32 => X"0621F562B1122DA70C3808458881056A5502AA150502828811FCD4EABDB1DFDF",
INIT_33 => X"96D55BBAAC55EAFAF86D35E4A92B4460D15060374FF72AAADF24559515705079",
INIT_34 => X"007FC0000007FC0000007FC07AAF12E00505D3FDF6A03D4BFB79AFA4C5CB5F58",
INIT_35 => X"0007FC0000007FC0000007FC0000007FC0000007FC0000007FC0000007FC0000",
INIT_36 => X"00000000000000000000000000000000000000007FC0000007FC0000007FC000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000040000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"212C001411984004084D000508C53810A03D1450E839B003342114428A000807",
INIT_01 => X"08000010400A0008010600000084004000400002000000000000000000140000",
INIT_02 => X"484DEBA0111800C004400D000000000028800001CC404E6008B4933336880010",
INIT_03 => X"CA1800080848B0423183089008C604224200000100A200002C280810098C0001",
INIT_04 => X"00000010822C00803804000001999EF9C00040B0002000001000640200001018",
INIT_05 => X"0000400244000000014200004000000004000000001000032000200002100800",
INIT_06 => X"208500000080412804100CB08000302220080408010000202000000404100844",
INIT_07 => X"5AF6FEF002230018010860C1833C460044204C000008A0041000080008202800",
INIT_08 => X"8D22C0F55000010000524481890BC000263000188AAAA10F8C1830562B25FC4C",
INIT_09 => X"B102002E20013600022D8819000000A000110A4000002C204000240420001000",
INIT_0A => X"02605C1C1108481200C000002040040820000020104100028800002801041001",
INIT_0B => X"081001004010810510040802040102008100200800A1100707040101E20BE0B0",
INIT_0C => X"58000003C0F000A000C4000003C0F000A000C0000012187087010AE4B0000000",
INIT_0D => X"04000003C0F000A000C4000003C0F000A000CC4200002F08E03080000010F180",
INIT_0E => X"0000000AAC00680000001F10E038000000078808C00000023461C0E000000127",
INIT_0F => X"5200040A00D000000202090C281F201803000000240218C0044200001E187806",
INIT_10 => X"400012900001EC03F000000000392100B00048230C200009A000130320480002",
INIT_11 => X"308000000961002880204A901C0E00000002C9000260640900004D0000904618",
INIT_12 => X"5C0C0312A002000000083881002880025A0A3C020000002A8400B00007806070",
INIT_13 => X"04080830008010468220A00008D0000801046004308A18500002012800090428",
INIT_14 => X"0840280206089000004090110200000000001454000200828008081110084000",
INIT_15 => X"4191AC191AC191A4191A00C8560C8D2910000060901010401E13405111220000",
INIT_16 => X"0410028000100800140000002004103224002006406401918C191AC191A4191A",
INIT_17 => X"2008020080200802008020080200802008020080200802008020080200800041",
INIT_18 => X"0080200802008020080200802008020080200802008020080200802008020080",
INIT_19 => X"0000000000000200802008020080200802008020080200802008020080200802",
INIT_1A => X"2431A589945201924924B060D757DF8A94102E038728287452B4008A04000000",
INIT_1B => X"75BADD6EAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8A28A28A28A28AB20",
INIT_1C => X"974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D2E974BA5D6EB75BADD6EB",
INIT_1D => X"00000000000000000000000000000000000303FFFFFFFFFFFFFFC00000BA5D2E",
INIT_1E => X"FDFFFA2FFD74000855555FFFFFFC01FF087BE8BFF5D2AAAB5555554000000000",
INIT_1F => X"EBFF455D04175FF5D7FEAAAA002ABDEAA5D2EBFFEFA2D17DEBAF7D1574BAAAFB",
INIT_20 => X"8415400005540155F7D16AB45002EA8ABA005540145557BFDEAA5500154AAAAA",
INIT_21 => X"5003DE00A2FFFFFEFAAD57DE00082AAAA00082A820BAAAD540145F7D5574BAAA",
INIT_22 => X"F7D5554AA5D2ABDEBA082A821455D2EA8B455D2A975EFF7AEBFF550055555FF5",
INIT_23 => X"FFF84155FFFFFFFFF55AAAABFFFF5D556AB45A2D16AABAAAAEBFE10AAFBD7545",
INIT_24 => X"10FF84174BA552EBDEBA0004020AA5D04155FFAAFFEABEFA2FBEAB455D7BD55F",
INIT_25 => X"F47015A800000000000000000000000000000000000000000000175FFF7D1400",
INIT_26 => X"FEAAF7D5524AAA2F0BAF7FABDFC7E10005F525D74BFBC51FF1471E8BEF55242F",
INIT_27 => X"50492490E17EAAA2AAB8F4515043DFC75575C7000B6AEBAEAA5D2EBDFFFBED17",
INIT_28 => X"B6FB6DF7DFD5038ABA140A2D00554517DEBDB6FB55142A8708202FBD257F1C75",
INIT_29 => X"AABFF55BC5B555C74B8A38E38085BE8B47A3A00503D1420AD000B420820AAE2D",
INIT_2A => X"AABD21EF1C2FEA5FDEBDB505FA4920AFE10082E925555F8FFDE38087FC51C7F7",
INIT_2B => X"1EFBFDBFF5FF1C00BF5D25475C7B7FEAFF45BEAABA4AF555168B68FEDF6AB52A",
INIT_2C => X"00000151EAE3D542A004380124921D20BFFFA0AA17AEB8BFF155552B6F5E8BFF",
INIT_2D => X"FF55516ABEFDD003EFE5093DC000000000000000000000000000000000000000",
INIT_2E => X"2BA5D2ABDFFFF7D57DEAAFFD5420B2A2D37DB07A3D795000087BC01458AFBC11",
INIT_2F => X"D608897FD610D01151C610592A974BAFBAC28B55550434D555C53E0CE2AAA874",
INIT_30 => X"3FE102400144ABAAFFF7DE772FDD56588042F72EF0851575FFAAFBDD5542B2ED",
INIT_31 => X"F6A81A239501755F504BDF557D79431FD006EABA100F3D68FFFAABAC20EF0400",
INIT_32 => X"55EAF57FF957CAAA7FABF7DFD0C6A7DFFFA07FC04EA0006BFE007E2E8315DD02",
INIT_33 => X"FADF6900FFFF68BEFDFFB4B1FE5551141E78A02803158517BD745AEAEA8FAF0C",
INIT_34 => X"0000000000000000000000165BAFBD542000D382964A92B403EE18D5408A6F2A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000040000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10E006600180111284380310006289800480032283E000A34301002001A0812",
INIT_01 => X"A145A00810790848048044A54E404340404000720885800802000906E4910200",
INIT_02 => X"5C010802020408040C455850AA055254090541A111200A104A0000000908B510",
INIT_03 => X"182002200C00004485264A001214912802150020218808002440854288890550",
INIT_04 => X"210302008014100120806B08702010102722C9E0412200651102418214049492",
INIT_05 => X"48416A98042912208552102442884882A58A08011290A1120A81230240018DCA",
INIT_06 => X"12800554528021C8023A28000031240048000100001170000155414109102066",
INIT_07 => X"000022104040810089080810211A04480420420154800088096A0EA8C0222080",
INIT_08 => X"080198C105424705510A08828A0B19080428040080A0A10F8102049300000804",
INIT_09 => X"3165541CD54822160A89E89020AA8AC4CA1D39CE215264B04040002400B80688",
INIT_0A => X"280201840548C80001C568146000001012D40D7182411080153801004800B057",
INIT_0B => X"4812050000080114100206000100818100900640C04C20104101021C00000310",
INIT_0C => X"00A00000010000A01001400000010000A0100801407234E34C1A980001552055",
INIT_0D => X"01400000010000A01000A00000010000A0100038000000000800000000405000",
INIT_0E => X"00000040A00002600000000010000000004608000850000000080000000001A0",
INIT_0F => X"400020C4000200420040000000001000000000002408000000A1000000020000",
INIT_10 => X"00001A04940000000000000020012800018000000000000D0288000000000003",
INIT_11 => X"0000000021480000508000000000000000400951000000000000681300000000",
INIT_12 => X"00000000000000000008600800004C000000000000000082A000015000000000",
INIT_13 => X"80004012C06000018004342AA000700000000000044000500000000022101800",
INIT_14 => X"958100134200904487400010022005E0110D524029263100009200151409130A",
INIT_15 => X"C9013C9011C90134901144801A4808AD4451394CD0391A541593C04B59084008",
INIT_16 => X"010400A0A890684444240120C0071420344423040240450114901149013C9011",
INIT_17 => X"080601806018060180200802008020080601806018060180200802048026C000",
INIT_18 => X"8000080001804018040180400800008000080601806018060180200802008020",
INIT_19 => X"1F83F03F03F00180401804018040080000800008000180401804018040080000",
INIT_1A => X"E90C042CB002102CB2CB2EE00271AE180616A85246C77250C7D00022012F81F8",
INIT_1B => X"28944A2504104104104104104104104104104104104104104104104104104608",
INIT_1C => X"128944A25128944A25128944A25128944A25128944A25128944A25128944A251",
INIT_1D => X"000000000000000000000000000000000003C3007FFFFFFFFFFFCE3F00944A25",
INIT_1E => X"EAA1055042AA105555421EFFFD568AAA002EBFEBA550002000AA800000000000",
INIT_1F => X"AA8BEFAAAE975FFA2D5555450851574000851554BAFFAE801FF087BE8BFF5D7B",
INIT_20 => X"2EA8AAA5D2EBFFFFA2D1554BAF7D17FEBAAAFFFDFFFA2D57DE10557BE8ABAF7A",
INIT_21 => X"D04175FFFFD5574AAAAAA974BA082EA8BEFAAD555555F7D568ABAF7D5574BA55",
INIT_22 => X"085557410F7AA97410087BD55FF087FEAA10A2FFEAAAA552AAAAAAAAAABFF455",
INIT_23 => X"05D7FE8B45F7FBFDE00085540155F7D56AA00007FEAA000055401555D7BFFE10",
INIT_24 => X"00082A820BAAAD540145F7D557410AA8428A10550017400550402155A2803FE0",
INIT_25 => X"000E28A80000000000000000000000000000000000000000000017400082AAAA",
INIT_26 => X"01FF1471E8BEF5574AFA00010ABFA38555F401D74BD16FAAA002ABFEAA550E82",
INIT_27 => X"FF400417FEF082F7AAA8BEFE2AA955EFA2DB5757FEAFBD2410005F57482E3AA8",
INIT_28 => X"F6DA82F7DF520385D2FE80AA5D2EBDFD7BED1574AAF7D5524AAA2F1FAF7FABFB",
INIT_29 => X"24ADAAAB6AAB8F455784155C75575C7000B6AE95492082EADBFFBEDB55555E3D",
INIT_2A => X"051C05571474024A81C5557578EBA087400007FC21C7005B6FB47F7A438E925D",
INIT_2B => X"E10A001FFB40038F68F7F578F7FFEF568E2808554717DEBDB6FA3D0075EDA800",
INIT_2C => X"000001043D1420AD000B420820AAE2DB4716DF7DFFDE381D716FA15550015428",
INIT_2D => X"AA002ABDEAA552A80010AAA88000000000000000000000000000000000000000",
INIT_2E => X"800087BD5410AAAA801FF55556ABEF5D517EEE00828FDEBA5D7BC015582D57DE",
INIT_2F => X"A2B2A3D169B07A3D7BFE10597BFDE00AEAC28BFFAAAE955EFAAFBC15F5A3D7D6",
INIT_30 => X"BDFEFFFFBC1154AAFFFFE107FF9D72A20842080BA5D2ABDF55F7D575EAAFFD50",
INIT_31 => X"97CF4780286A2105D2A3FEBAFFAC28B555504145555A53C00B2A2AA02000082A",
INIT_32 => X"FFFDA02003FFDEAA8557D65550915544AA5D51574EAA28015400547FC315D007",
INIT_33 => X"16F9E2555500174AA282E20BFFFF842AAAAADD5699ADABD5A8AAA0051575FFA2",
INIT_34 => X"0000000000000000000000030EF04003FE102400144ABAAFFD75E7F2BDDD2B80",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000080000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"210C44A20020248B08431120001604B8156023104C4077133420400A02380202",
INIT_01 => X"200C9A424080216D3C2462C99E104B49404040028804A0080A000416A8D90A0C",
INIT_02 => X"4809A902031800444461089C66E331352180D468B8240E600C0081110B80ACD0",
INIT_03 => X"DA16C2210C0001D231A30A0648C68428320066010A80881068A80C401CC46330",
INIT_04 => X"2088601DA82700EC92307064A3756910088469A01C250210990240420E005A48",
INIT_05 => X"2D2060182414411A314A0A02C18C01B9854368080A506912018C2502484038D1",
INIT_06 => X"16801CCCAA8061E8061C0D008020140520080769000420202133CCC50C110804",
INIT_07 => X"5800B65040630008810C20508138071604A461833280038C89904E6400232008",
INIT_08 => X"0800906010521D1CC80204918949540C061000088000A90F840A50963A017845",
INIT_09 => X"A037A02C68552A35620C88900A69876100810A6A84C82C400040300D40D20A48",
INIT_0A => X"062A10B40042C80000CCE4CC2045051913208CE80243048008204100402079CC",
INIT_0B => X"C81301004C18912102060C0207010201C190200400A401042D00F15884030170",
INIT_0C => X"0190148000000800100450148000000800100401CB33494594532980733322CC",
INIT_0D => X"05101480000008001004F014800000080010051C000040000000000000480000",
INIT_0E => X"00000044000001680180400000000000014000000B1004090000000000040080",
INIT_0F => X"00812E44000024400140800280000000000002000008000001B0000040000000",
INIT_10 => X"0002080CCC0002000000000020401000034010480000010402D8040440000041",
INIT_11 => X"00000000601000064180104400000000004100570080880000082015C0209000",
INIT_12 => X"00820080000000000100401000061C0001000000000000904000094C00201800",
INIT_13 => X"4408400000A26285A03224E670094008010000004444010E2050000420801880",
INIT_14 => X"4DC10283429294408740C0B48202854C011CD75C0102A30400A8891451284B26",
INIT_15 => X"4901A4901849018C901A648056480C2D4449116DC0115C41159B655F112AC008",
INIT_16 => X"0510000000DA690C1D20030BA0011421B404220402404501A49018490184901A",
INIT_17 => X"280803808038080380803808038080380C0280C0280C0280C0280C0680C28051",
INIT_18 => X"00C0280E030080380A030080380A030080380C0280C0280C0280C0280C0280C0",
INIT_19 => X"B556AA9556AA830080380A030080380A030080380A0200C0280E0200C0280E02",
INIT_1A => X"742C000A981E80249249206018F18E0C85142822266800586291000A844D54AA",
INIT_1B => X"A9D4EA7524924924924924924924924924924924924924904104104104104A20",
INIT_1C => X"1A8D46A351A8D46A351A8D46A351A8D46A351A8D46A351A8D46A753A9D4EA753",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF849010D46A35",
INIT_1E => X"42000AA802AA10F7D57FEAA557BE8B45A2D5555EFAA800015508000000000000",
INIT_1F => X"BC0155A280021EFA2FFE8B4555042AA105555421EFFFD568AAA002EBFEBA5551",
INIT_20 => X"D5574000851554AAFFAE801FF087BC01FF5D7FEAA10550402000AAD56AAAA557",
INIT_21 => X"AAE975FF005540145A2D157410AAD17DFFF5D0400010AA842AAAAFFD542000FF",
INIT_22 => X"F7AE975FF080428B455D7FFDEAA5D55574BA00517DE105551420BAF7AAA8BEFA",
INIT_23 => X"F007FFFEAAAAD5554AA552EBFFFFA2D5554BAF7803DEBAAAFFFDFEFAAD57DEAA",
INIT_24 => X"EFAAD555555F7D568ABAF7D5574BA552E800BAAAAE800AA087BD5555552A821E",
INIT_25 => X"155080E800000000000000000000000000000000000000000000020BA082EA8B",
INIT_26 => X"FAAA002ABFEAA555E02000E28AA8A38EBD578E82E975EAB6DBEDF575FFAA8E02",
INIT_27 => X"87A38AAD56DA824975C217DAA84021FFAAF5EAB55EBAEADA38555F451D7EBD16",
INIT_28 => X"E2DABAFFDB47412ABFE90410005F57482E3AA801FF1471E8BEF5575EFA00012A",
INIT_29 => X"5F47082E3AAA8BEFA02A955EFA2DB5757FEAFBD2400BED57FFD7410E05038BE8",
INIT_2A => X"2F1FAF7FABFBEAE2AEBA4974871C043AB6D4975FFEBA5D71D742A407FFFE0055",
INIT_2B => X"1C75D25C74920821D708757AE2AA3FFC04AA552EBFFD7BED157482F7803AEAAA",
INIT_2C => X"0000007092082EADBFFBEDB55555E3DF6DA82F7DF7AE38497FC00BAB6A485082",
INIT_2D => X"FFFFFFD75FFAAAE8014500288000000000000000000000000000000000000000",
INIT_2E => X"EBA5D7BD5545A2D57DEAA002EBDEAA557BC0010AAA8A8ABAAAD568A1020516AB",
INIT_2F => X"29EF5C517EEE00828D74AAFBD57DE000057C21FFAA80001FFAAD57EB55A2A8AB",
INIT_30 => X"7DF55082E974AAFFAABDEBA77FDD66A0ABBDC2000087BD5410AAAA801FF55556",
INIT_31 => X"7C14100957FF6105D7BD5400AAAC28BFFAAAE955EFA8FBC15E5A3D5D7400FFD5",
INIT_32 => X"D1554A8FFC42AA10A7D169F57ABD7FEEBAAA841550555002ABFF54517EEB25D5",
INIT_33 => X"96F014AAFF84154105555C215500000014558557FA42A3D7020BA5D2ABDF55F7",
INIT_34 => X"000000000000000000000015400082ABDFEFFFFBC1154AAFFFFE10FFF9DF2020",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000040000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A108400020612C80284210081034849800A000303100048B3432C82904204002",
INIT_01 => X"010398000008004C1C20650E1E104348403008418984014902030006A0910200",
INIT_02 => X"480108A200000000444048E41E80F00A4104311868200200080000000988A390",
INIT_03 => X"0CA08220080000D004060A0240101028270012603000000030808C0208C000F0",
INIT_04 => X"4403A609A055306BC2C0735810CEE5100A0A40E06B8360E3808241D03845D002",
INIT_05 => X"ECE0498800791403AD3038AE079059A790E245819A41E4120BAB87800001D312",
INIT_06 => X"06000C3D220003E0001A210088B1008C4004034912120000010FC3C00000A064",
INIT_07 => X"5000220440000000090800002118400204206100F040018019004B8001232088",
INIT_08 => X"0810884441123323C0424180880B0108002000000880890F9000041200000845",
INIT_09 => X"230B6715A4786E0F5A8C889031EF9F45D884794FA03A24781840100D000E1140",
INIT_0A => X"0C4202200142400004DC3C82600401003200872003FB1400082840001022003C",
INIT_0B => X"C800940008088034040000010000808140901000C00001008800A01814000840",
INIT_0C => X"02E0100000000800000620100000000800000001C07261841840310240F070C3",
INIT_0D => X"0680100000000800000760100000000800000435100040000000000000080000",
INIT_0E => X"00000004000000D8008000000000000001000000155000080000000000040000",
INIT_0F => X"000100EC00004002214000008000000000000200000000000094100040000000",
INIT_10 => X"000200010C000200000000000040080005800008000001000368000040000040",
INIT_11 => X"000000004008000448000040000000000001007C000008000008001D00001000",
INIT_12 => X"000000800000000001000008000017000100000000000010200002C800000800",
INIT_13 => X"0000549000027200800E271E00288400800208004804C0080000000052800800",
INIT_14 => X"454000924280D144B14041340A880EC51160525C0022510006BE1002C6150F5E",
INIT_15 => X"010C1010C1010C3010C14086980861AD447F2201D899BA403593514B59A30088",
INIT_16 => X"010448002098694C15204369E00116203445E3443043410C5010C3010C1010C3",
INIT_17 => X"180000006018000000200804010020080400002018040000600800010064E000",
INIT_18 => X"8060000001000008060180201000000040180001006008000100201804000020",
INIT_19 => X"934D964C32698000401802008060000401000008060080201004000000080201",
INIT_1A => X"0991A185145019A28A289830C700FC0A0002870BB5ED0B34504048828464B261",
INIT_1B => X"351A8D46AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8A28A28A28A28AF4C",
INIT_1C => X"8341A0D068341A0D068341A0D068341A0D068341A0D068341A0D46A351A8D46A",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8EE3EC1A0D06",
INIT_1E => X"40155080000155FF843FFEFAA84001FF5D043FEAA5D55420AA002A8000000000",
INIT_1F => X"A80010FFAE975FFAA80001EFA2AAAAA10F7D57FEAA557BE8B45A2D5555EFAAD1",
INIT_20 => X"AAAAA105555421EFFFD568AAA002EBFEBA555542000AA80001555D04174AA002",
INIT_21 => X"280021EFA2FFE8B45F78400145FF842AAAAA2AA800BA5D51555EF002AA8BFFAA",
INIT_22 => X"00003DFEF080428B455D002AABA5D2AAAAAA5D2E82000AAD568AAA557BC0155A",
INIT_23 => X"FAAAAA8BEF552E820000851554AAFFAA801FF087BC01FF5D7FEAA105D0428B45",
INIT_24 => X"FF5D0400010AA842AAAAFFD542000FFD57DF55A280154BAA2FBE8AAAF7AA821E",
INIT_25 => X"092142E00000000000000000000000000000000000000000000015410AAD17DF",
INIT_26 => X"AB6DBEDF575FFAADE02155080E85145E3803FFEFA284051D755003DE92415F42",
INIT_27 => X"851455D0A124BA002080010FFA4955C7BE8E021C71C0A28A38EBD57DE824975E",
INIT_28 => X"B505D71424AABD7F68E2FA38555F451D7EBD16FAAA002ABFEAA555F42000E2AA",
INIT_29 => X"D56DA824975C217DAA84021FFAAF5EAB55EBAE82145F7802AABAA2A480092415",
INIT_2A => X"575EFA00012ABFB6D080A3AFEF080A2FB45490E2AA824924AAA92550A07038BE",
INIT_2B => X"AAFFEAA00F7AE821D7B6A02FBC71D0E10010005F55482E3AA801FF1471C01EF5",
INIT_2C => X"0000010400BED57FFD7410E05038BE8E2DABAFFDB6FA12ABAEBDF7DAA80104BA",
INIT_2D => X"4555043FE10087BC2000552C8000000000000000000000000000000000000000",
INIT_2E => X"ABAAAD57DE1000516ABFFFFFBD75FFAAFFC0145002897555A2803FFFFAA84175",
INIT_2F => X"DEAA557BC0010AAA895555042E820BA080400010FF8017545F7AE821455D2CAA",
INIT_30 => X"2AAAAAA8002010007FC0155D5022A955FFACBFEBA5D7BD5545A2D57DEAA002EB",
INIT_31 => X"43CAB0552C97CAAFFD57DE000057C21FFAA80001FFAAD57EB55A2A880155F780",
INIT_32 => X"AA801FF5555421EF58517EAB00028A9BEF002EAABEF002EBDF45542AAAA00080",
INIT_33 => X"A90FDFEFA280020BAA2FFEAA10FFAE82145F7803CFE55D2CC2000087BD5410AA",
INIT_34 => X"000000000000000000000002000FFD57DF55082E974AAFFAABDEBAF7FDDE6A0A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000080000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50DF4A0791B3FCB694379283C81FD996A091832102004A337A20E07C0C1E006",
INIT_01 => X"295FBC448000804C5C6A60000C34C26841280A00084000C8C212802EE2953235",
INIT_02 => X"C809AD5EB118E640A4D158FC011FF0002080000082E8C66609DB7DDDCB1FA036",
INIT_03 => X"4A120E4C3A4C90D214A35E824852857A0A20640A88800000B8E0FC52A884500E",
INIT_04 => X"001440809A2604005934800041110A71E290E8B010DB221C662AE22DC0AA3448",
INIT_05 => X"12026A2A1B88C31841CDC451B860A6507BEBD18A65AE10571450DE8112522449",
INIT_06 => X"80752C03736281D628398CD0A4C894EA2054237F271331095100D82D0C2C82A2",
INIT_07 => X"5E64B66BD6231CC81529A356AD3AC601C57FF54FF149A46490261C4B39203F70",
INIT_08 => X"AD0099410015814FC602C4B1B93947F8621030C800001D7FA46A95172E937835",
INIT_09 => X"2C836D35B68D26C082DE9AB88C104020000208401807B78739010C04E17F5014",
INIT_0A => X"082099129008F25615C3FC01A2102109204C28B6706168128920C469E7C00A00",
INIT_0B => X"E92C23E210A0B246C2234010A108D0042811461C0401502644A40106C14FD22A",
INIT_0C => X"E00BF1BFE1F000BE1FC40BF1BFE1F000BE1FC80028120800800100653FF0313F",
INIT_0D => X"040BF53FE1F000BE1FC40BF53FE1F000BE1FCC806FFFEF0AE83080E2AEF2F1F1",
INIT_0E => X"013879FAAF8FC003FEDF5F12F0380231F0FF963F00A7FBDF3669C0E008C3CBFF",
INIT_0F => X"F2008022CBAC8B9DDEB779BEA91F30180309A0F83FEAB8FC7C006FFFDF1A7806",
INIT_10 => X"4131BF940DFFFE03F00003F03FB929E9C19BE8EB0C2098DFE2EF7B2760483137",
INIT_11 => X"3080E29F3B69E9F4427EEED41C0E004C72FEC95DEFE46C090626FF1537F15618",
INIT_12 => X"FC0E0392A0024B83F07F7989E9F01DFFFB0A3C0202B877EAA7A7C1CBFFD07870",
INIT_13 => X"C0404020040001C4E7F1787E0C8028514885C566241902508C83A7D1B7EFAC6D",
INIT_14 => X"4DF46A170F92C7E20F0430938008AC38C4184B100136858C9298A8560688F4C1",
INIT_15 => X"6B8C86B8CE6B8CA6B8CC15C6435C670C10EB4124D2B3903BF5C9710C1191DCA0",
INIT_16 => X"2030461200984D041C40208400230E71B3104E5636E3178C86B8CC6B8CA6B8CE",
INIT_17 => X"0040118401184610042110401184410846110421104010844118421504238200",
INIT_18 => X"8441184011844100461004211046100461084211042100441084011842100461",
INIT_19 => X"DA6924965B4D1004610840118401084410840110421004610046110421084410",
INIT_1A => X"FF9FBFAF2DDA3B9E79E7BED9CFEF73B6FFE74FC3F78FFF6DB7ED438A183124B2",
INIT_1B => X"DDEEF77BBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEDFD",
INIT_1C => X"BDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BBDDEEF77BB",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF853FB5EEF77B",
INIT_1E => X"020AA002AAAABA555140155087FFFFEF00042AB555D2E955FFF7FFC000000000",
INIT_1F => X"E975FF5D5568B555D7BD5545FFD540155FF843FFEFAA84001FF5D043FEAA5D04",
INIT_20 => X"FFEAA10F7D57FEAA557BE8B45A2D5555EFAAD5401550800001FF5D00001555D2",
INIT_21 => X"FAE975FFAA80001EF002AAAABAF7D168A10A2D17FF45A2FFC0000AAAE974AAFF",
INIT_22 => X"F7803DF55FFAEBFE005D2EAAB45557BD55555555401555D04174AA002A80010F",
INIT_23 => X"5552E955EF5D7FEAA105555421EFFFD568AAA002EBFEBA555542000A28028BFF",
INIT_24 => X"AAA2AA800BA5D51555EF002AA8BFFAAAA820AA5D517DF55082E974BA087FE8B5",
INIT_25 => X"5C7F7FBC0000000000000000000000000000000000000000000000145FF842AA",
INIT_26 => X"51D755003DE92410F42092142E28ABA5D5B4516D007FFFFFF1C042FB7D492A95",
INIT_27 => X"851C75D0E02145492E955C75D5F6DB55497BD5545E3DB45145E3803AFEFA2840",
INIT_28 => X"BC7028A2AA95492FFFFE8A38EBD57DE824975EAB6DBEDF575FFAADF42155082E",
INIT_29 => X"0A124BA002080010FFA4955C7BE8E021C71C0A2DABAF7D16DA28A2DB7AF7DB6F",
INIT_2A => X"55F42000E2AAA8BEFE3843AF55E3AABFE105520AFB45557BD5555415F4514549",
INIT_2B => X"082E954AA087FEDB7D5D2A155D7157BEFA38555F451D7EBD16FAAA002ABFEAA5",
INIT_2C => X"0000002145F7802AABAA2A480092415B505D71424821D7F68E07082495B7FF7D",
INIT_2D => X"EF5D003DFEF002E95555F7FDC000000000000000000000000000000000000000",
INIT_2E => X"555A2802ABFFAA841754555043FE10082A82000552CAAAAA5D7FD75EF087BFDF",
INIT_2F => X"75FFAAFFC0145002895545552E80145002E955455D7BFDF45007FD7555A2F9D5",
INIT_30 => X"7FEAAAAFFEABFFF7FFD54BAA2AA95410F7FDEAABAAAD57DE1000516ABFFFFFBD",
INIT_31 => X"BD55550879D5555002E820BA080400010FF8017545F7AE821455D2CBFEAAFFD1",
INIT_32 => X"D57DEAA002EBDEAA557BC0000AAA8A8BEFA28028B45AAAABFE0009043FF555D7",
INIT_33 => X"FAC97400087FFFFFF002E954AA087BFFFFF5D2E975455D7DFFEBA5D7BD5545A2",
INIT_34 => X"000000000000000000000000155F7802AAAAAA8002010007FC0155550222955F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000300000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B0061A258A2840112C03002C180004003220200403302301C0381A0082",
INIT_01 => X"860041C838394848008100000042026041000000090800090210010000510204",
INIT_02 => X"080108220C1000004464080000C008010000000001243240080080000988A050",
INIT_03 => X"080000010C23404080020A600200002983800504488000103080050C08C10000",
INIT_04 => X"0040504280A682104011230010000010002040E9102050101000400A00003000",
INIT_05 => X"0409400984008000414A00014000002004100020005004020010204044802800",
INIT_06 => X"301223FC028911E8911900000224200248A653E908C0248489FF000809108000",
INIT_07 => X"0000220441820000090C080001184400142040200E824008900008000220600A",
INIT_08 => X"1A18946451007FA0380200808809010C182000000000090F8100001220000804",
INIT_09 => X"300240B4A409223F020988100808200490142B441BF82C20401481540A000008",
INIT_0A => X"264285180542408000D001BE090693912000002004410489080001100017E2FD",
INIT_0B => X"091081090A4491A40052A129519428CA142288010A5A21214601F01A220602A0",
INIT_0C => X"18100400000000A00034100400000000A00033A00813004104020818800F2400",
INIT_0D => X"F4100080000000A00034100080000000A0003142000000000000000000055D00",
INIT_0E => X"00000001E8002900010000000000000000066000C20004000000000000000120",
INIT_0F => X"4D240C2000502000000080000000000000000000240146800142000000000000",
INIT_10 => X"00001260F0000000000000000007F00032201000000000091A00040000000002",
INIT_11 => X"0000000005D00008958010000000000000003F4000008000000048D240008000",
INIT_12 => X"008000000000000000082670000CC0000000000000000007C000301400200000",
INIT_13 => X"0120849A5250101482202301F05101202420000810C219500150002800101280",
INIT_14 => X"454110030212C140011204D020880C000018431DE802015022A62A1596C8B580",
INIT_15 => X"016C2016C2016C6016C440B6000B600C446B0104D09192013589701C59800002",
INIT_16 => X"51804A0028904C425016040820978221B0000005B05B416C0016C0016C4016C4",
INIT_17 => X"8CA3294A528CA328CA1294A528CA3284A5294A728CA3284A529CA728CA100508",
INIT_18 => X"CA3284A129CA7294A328CA1294A729CA128CA329CA5294A128CA3294A5294A32",
INIT_19 => X"1C71C718638E28CA529CA7284A128CA7294A528CA1284A729CA1284A3284A529",
INIT_1A => X"ED9DBDAFBC5E9BBEFBEFBEF9CFF1FE1E9F52AFF9F3E77B7CF7F40A00107638C3",
INIT_1B => X"FCFE7F3F8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E76C",
INIT_1C => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9",
INIT_1D => X"00000000000000000000000000000000000303007FFFFFFFFFFFC61AC8FE7F3F",
INIT_1E => X"955FFF7FFC21EFF7D17DEAA5D2AAAAAA5D557DE105D2EBDF55557FC000000000",
INIT_1F => X"03DEAA5D5568BEF5D042AA10A2AAAAABA555140155087FFFFEF00042AB555D2E",
INIT_20 => X"5540155FF843FFEFAA84001FF5D043FEAA5D00020AA002A82145555542010FF8",
INIT_21 => X"D5568B555D7BD5545FFD568AAA5D00154AAAAD1420BA00557DF455D7BFFEAA55",
INIT_22 => X"F7843FF55007FFDEAAA284020BAAAD168BFF0800001FF5D00001555D2E975FF5",
INIT_23 => X"5AAAEBFE10FFFFEAA10F7D57FEAA557BE8B45A2D5555EFAAD540155080000000",
INIT_24 => X"10A2D17FF45A2FFC0000AAAE974AAFFFFC21EF5551401EFF7842AA00FF841754",
INIT_25 => X"F45497FC000000000000000000000000000000000000000000002AABAF7D168A",
INIT_26 => X"FFFF1C042FB7D492A955C7F7FBC71EFFFD57FE825520ADA92495B7AE10412EBF",
INIT_27 => X"0716D415F47000F78A3DE92415F6ABD7490A28A10AAAAA8ABA5D5B4516D007FF",
INIT_28 => X"F78F7D497FFFE925D5B45145E3803AFEFA284051D755003DE92410E02092140E",
INIT_29 => X"0E02145492E955C75D5F6DB55497BD5545E3DB6AA92550A104AABED1470AA005",
INIT_2A => X"ADF42155082E87038FF8038F6D1C7BF8EAAAA80020BAA2DB68BC7140E051C75D",
INIT_2B => X"FF8428A00E38412545AAAE3FE10A3FBE8A38EBD57DE824975EAB6DBEDF575FFA",
INIT_2C => X"000002DABAF7D16DA28A2DB7AF7DB6FBC7028A2AA95492FFFFC71EF415F471C7",
INIT_2D => X"00007FEAA10002ABFF450079C000000000000000000000000000000000000000",
INIT_2E => X"AAA5D7FD75EF087BFDFEF5D003DFEF002E95555F7FDD55EFF7D57DE005D003DE",
INIT_2F => X"FE10082A82000552C955FF007BD5410FFAABFE00087BE8B45082EAAA10A2A8AA",
INIT_30 => X"820AAF7D5574AA087BEABEF007FFDE00557DD5555A2802ABFFAA841754555043",
INIT_31 => X"BEAB55552C95545552E80145002E955455D7BFDF45007FD7555A2F9EAA005D2A",
INIT_32 => X"516ABFFFFFBD75FFAAFFC01450028974BAFF842ABFF557BE8ABAA284020BAA2F",
INIT_33 => X"7FDD55EF007BD5555F7802AA10AA8000145AAAEBFE10A2F9EAABAAAD57DE1000",
INIT_34 => X"00000000000000000000003FEAAFFD17FEAAAAFFEABFFF7FFD54BAA2AA95410F",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000240000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10844B00482258A2842112C024504188000003000000003302300C018180006",
INIT_01 => X"020008422008604D042080000211024840000000080000080200080000110204",
INIT_02 => X"4801082048100000444008040080000041000000000222400800000009000010",
INIT_03 => X"0802030288A148D0000208424000002103006400088000003080000408C10000",
INIT_04 => X"00004000890600004032030010000010008060E4100000140006500800403040",
INIT_05 => X"0400400080000018414800810000002000000000004000328010000080882000",
INIT_06 => X"281A8001220021E0021803000224200200000360888420000000100808000000",
INIT_07 => X"5000220409020000090800000118040014A061200052500810000C490323208E",
INIT_08 => X"1A9098411110014000424090980B0002102000000000010F8000001220000805",
INIT_09 => X"31024034A4092200820D899408000004D0143B4410002C800080020450800001",
INIT_0A => X"24028011444240A88CC00100200D0010200008B2066397014800221400140C01",
INIT_0B => X"080001000C008124000000000100008000100404204C25200451A01A00A620A5",
INIT_0C => X"1C0014800000F001E02C0014800000F001E021141213000000000010B0001000",
INIT_0D => X"CC0014800000F001E02C0014800000F001E022420000400004C3201C51040908",
INIT_0E => X"60078601084038000180400002C0E00E0E004100E000040900000B0380383400",
INIT_0F => X"08146800105100000000800284004160C0301D07001504820242000040000198",
INIT_10 => X"908C404AFC000200030F000FC00610103BE0104810C8462014F8040446120C88",
INIT_11 => X"C3201C608410100FD5801044013098038D00309F008088C2419100A7C0209021",
INIT_12 => X"00B2048902C0807C0E008450100FDD000100411C8107880440403DDC00201804",
INIT_13 => X"00100496406010A0A2002200125140000000221110C018066250402E32901A80",
INIT_14 => X"454214028220141530400910CA800900326790500002001444001C0050140A00",
INIT_15 => X"5120551205512055120708901A8901A104804000801212541403C15178008010",
INIT_16 => X"01004200A09A49445420000DC000152804C9A384814809201512015120151201",
INIT_17 => X"0004000000080200806008020000000000000020080200802000000000008000",
INIT_18 => X"0000000000802008000000000002008020000400000000000080600802008000",
INIT_19 => X"0002082080000100000802008020100000000008020180000000000020180200",
INIT_1A => X"0000000000000000000000000000000000000000000000000005428A14584104",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8DD9EC000000",
INIT_1E => X"BDF55557FFDE00557BEAABAA2AEAABEFF78015555AA801741055554000000000",
INIT_1F => X"BEAAAAAAD157555AA803FEBA5555421EFF7D17DEAA5D2AAAAAA5D557DE105D2E",
INIT_20 => X"802AABA555140155087FFFFEF00042AB555D2E955FFF7FFD5555557BEABFFF7F",
INIT_21 => X"D5568BEF5D042AA10A2AA955EFF7FFD5400F7FFFDFEFAA80000BAAAAA820BAA2",
INIT_22 => X"5D7FE8A000004154BAF780001EFAAAAA8B45000002145555542010FF803DEAA5",
INIT_23 => X"5AAD5555EF557FC0155FF843FFEFAA84001FF5D043FEAA5D00020AA002ABDEBA",
INIT_24 => X"AAAAD1420BA00557DF455D7BFFEAA5555575455D2AAABFF5551421FFAAD15754",
INIT_25 => X"4385D5540000000000000000000000000000000000000000000028AAA5D00154",
INIT_26 => X"DA92495B7AE10412EBFF45497FFFE385D71E8AAAAAA0A8BC7EB8417555AA8410",
INIT_27 => X"D056D5D75EABC7FFF5EAAAABEDF5257DAA8438EBA4155471EFFFD57FE825520A",
INIT_28 => X"0070BAA2A0870BAAA8028ABA5D5B4516D007FFFFFF1C042FB7D492A955C7F7FB",
INIT_29 => X"5F47000F78A3DE92415F6ABD7490A28A10AAAA925EFEBFFD2400EBFBFAFEFAA8",
INIT_2A => X"10E02092140E3DE924171E8A281C0E10482F784001D7AAA0AFB6D1C040716D41",
INIT_2B => X"4955421EFA2DF5557DAAD5D05EF0175C5145E3803AFEFA284051D755003DE924",
INIT_2C => X"000002AA92550A104AABED1470AA005F78F7D497FFFE925D5B525454124AFBC7",
INIT_2D => X"55A28015545A284000BA5D534000000000000000000000000000000000000000",
INIT_2E => X"5EFF7D57DE005D003DE00007FEAA10002ABFF450079FFEAA5D5568ABAA2842AB",
INIT_2F => X"DFEF002E95555F7FDC01EF55556AB55F7D56AABAF7FBC01EFA2842AABA085755",
INIT_30 => X"C2000A2FFEABFFAA84174BAAA80174AAAA862AAAA5D7FD75EF087BFDFEF5D003",
INIT_31 => X"43DFEF5D02155FF007BD5410FFAABFE00087BE8B45082EAAA10A2A8801FFA2FF",
INIT_32 => X"841754555043FE10082A82000552CBFE10085168AAA552A80010F78000145AA8",
INIT_33 => X"57DC014500003FF450051401FFA2FBD55EFAAD5421FF085755555A2802ABFFAA",
INIT_34 => X"00000000000000000000002AA005D2A820AAF7D5574AA087BEABEF007FFDE005",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0000040042840002C00000018000002700500030B3132000400812082",
INIT_01 => X"A14008420008204D042100000212026840000000180800080200090048510200",
INIT_02 => X"080108020090000004655C000080000051000000002402400800000009008010",
INIT_03 => X"0002000100300C408422420002108108028065044880001030808D4288C10000",
INIT_04 => X"0002504688A28210003100000000001002A0E88910A032541000090A00643040",
INIT_05 => X"04092A081400D118410A002140004020140001A9005000004810A1C0044D2800",
INIT_06 => X"0010EFFD228931C8931820002080258A48A653E00213248C98FFC0094910A222",
INIT_07 => X"4000220440120000090C0810210A040034A040000046180810000C4907036008",
INIT_08 => X"50D88C2450000140004200808809000C012000000000010F8102041320000000",
INIT_09 => X"2002002020010200828C88020800200040801A40100228A1585481544A804040",
INIT_0A => X"A20804802400C80080D0010029069290200008B20E2304086800400640200801",
INIT_0B => X"091084090A4C81240251A328D094684B34A288050A5828012009504420102180",
INIT_0C => X"080004801E0FF00010000004801E0FF000100220021200000000000080001000",
INIT_0D => X"000004801E0FF00010000004801E0FF000100440000000F517CF600000400104",
INIT_0E => X"E000004008100800010040ED0FC7E000004008804000040109963F1F80000080",
INIT_0F => X"0020040020100000000882431660CFE7C0F00000000800810040000000E587F9",
INIT_10 => X"B0000808000001F80FFF0000200008021040134473D800040010045C1F360001",
INIT_11 => X"CF600000200802028001102EA3F1F80000400002008B83D6C0002000802688E7",
INIT_12 => X"03F2DC2D1FC18000000040080202800004D5C3FD80000080200818000027928F",
INIT_13 => X"0122C01A52501094222002000110012064200008848218002100100C00004112",
INIT_14 => X"4500048240C08400841204D0A00089000100001DE9248104300294428148A480",
INIT_15 => X"4800048000480004800004002240020850884000901210140011C010312B888A",
INIT_16 => X"51A4C000889A4D0E1D7624086491800420044240020004004480004800048000",
INIT_17 => X"84A1284A128CA328CA328CA328CA328CA328CA1284A1284A1284A12C4A14E508",
INIT_18 => X"CA328CA3284A1284A1284A1284A328CA328CA328CA328CA3284A1284A1284A12",
INIT_19 => X"000000000000284A128CA328CA328CA328CA3284A1284A1284A1284A328CA328",
INIT_1A => X"4799B1A014503EB65B6594F14A87D78AF421448BB528AF75D640088884400000",
INIT_1B => X"7C3E1F0F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79EDFC",
INIT_1C => X"87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F4F87D3E1F0F87C3E1F0F8",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF834FA53E1F4F",
INIT_1E => X"174105555420000000021EFAA843DE00F7803FEBAFFFFC2000557FC000000000",
INIT_1F => X"43DE005504175FF08514014555557DE00557BEAABAA2AEAABEFF78015555AA80",
INIT_20 => X"7FC21EFF7D17DEAA5D2AAAAAA5D557DE105D2EBDF55557FD54AAA2AA955FF000",
INIT_21 => X"AD157555AA803FEBA55556ABFFA280154BAFF803DF45FFD17DFFFFFD56AA0055",
INIT_22 => X"002AAAAAAA2D57DF450004154BA087BEAAAAF7D555555557BEABFFF7FBEAAAAA",
INIT_23 => X"5FFD1555EFA2802AABA555140155087FFFFEF00042AB555D2E955FFF7FFD5410",
INIT_24 => X"00F7FFFDFEFAA80000BAAAAA820BAA280000AAA2843DE1008556AA00A28028B5",
INIT_25 => X"0285D75C00000000000000000000000000000000000000000000155EFF7FFD54",
INIT_26 => X"8BC7EB8417555AA84104385D5542038000A001C7A2803AE38FF843DEBAEBFFC2",
INIT_27 => X"D24BAA2AA955C708003FE285D00155FF0055451555D5F7FE385D71E8AAAAAA0A",
INIT_28 => X"B78FFFE3DF6DA284175C71EFFFD57FE825520ADA92495B7AE10412EBFF45497F",
INIT_29 => X"75EABC7FFF5EAAAABEDF5257DAA8438EBA415568BEFA28E124AAF7843AF7DEBD",
INIT_2A => X"92A955C7F7FBD54380020ADA82BED57DF450804104920875EAA82F7DB5056D5D",
INIT_2B => X"005F68A10BE802DB55E3DB555FFF68028ABA5D5B4516D007FFFFFF1C042FB7D4",
INIT_2C => X"00000125EFEBFFD2400EBFBFAFEFAA80070BAA2A0870BAAA80070BAA2803DE00",
INIT_2D => X"AAFF803DEBAAAFBC20BA55514000000000000000000000000000000000000000",
INIT_2E => X"EAA5D5568ABAA2842AB55A28015545A284000BA5D53420BA082E82155AA802AA",
INIT_2F => X"AA10002ABFF450079C20BAAAAE9754500043DEBA5D04175EF0855575455D7BFF",
INIT_30 => X"820AAFF802ABEFAAFFEABEFAAFFFDEAA0051555EFF7D57DE005D003DE00007FE",
INIT_31 => X"16AA10FFFFC01EF55556AB55F7D56AABAF7FBC01EFA2842AABA085768BFFA2AE",
INIT_32 => X"7BFDFEF5D003DFEF002E95555F7FDD74BA08043DE10F7D17FF55000000010085",
INIT_33 => X"A86174AAAA843DE00087FE8A00F7843FF45AAFFD75EFF7842AAAA5D7FD75EF08",
INIT_34 => X"0000000000000000000000001FFA2FFC2000A2FFEABFFAA84174BAAA80174AAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000100000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000B0001800002840002C0000281800000030000000033022000000000006",
INIT_01 => X"000009801830084C182060000C104268413C0A61590001D90213C00000110200",
INIT_02 => X"680108200010000054400C000080000041000000010002400800800009082011",
INIT_03 => X"0008000004002040000200100000000042800584488000103081880008800000",
INIT_04 => X"00005842802AC210001000000800001000004080100040140080040800003100",
INIT_05 => X"0400000040000080410800010001002000000000004000002010000040002000",
INIT_06 => X"10100001221911E1911902000020200201A2D3E8000C2C84880010080800004C",
INIT_07 => X"C0002204000200000B080000010C040004A0400000C0000810000C5901036000",
INIT_08 => X"002A84300000014000C2008088090000002000000000030F8000001220000408",
INIT_09 => X"210000020000120082088801080020400000084010002880000C803400000008",
INIT_0A => X"020000040000480100D0010019019190200008B2022380800802010000000801",
INIT_0B => X"09000119064C810500D0A36851B428DA14368C801A1400000100500400000090",
INIT_0C => X"08100080000000A00000100080000000A00000000212000000000000B0001000",
INIT_0D => X"00100400000000A00000100400000000A0000540000000000000000000005100",
INIT_0E => X"00000000A8000900000040000000000000060000420000010000000000000120",
INIT_0F => X"4000040000102000000000020000000000000000240000800140000000000000",
INIT_10 => X"00001204FC000000000000000001280013A000400000000900E8000400000002",
INIT_11 => X"0000000001480004D5800004000000000000091D008000000000480740200000",
INIT_12 => X"0002000000000000000820080004DD000000000000000002A00011DC00001000",
INIT_13 => X"0322C01032301006022082000010032024200000048019500000000832901A80",
INIT_14 => X"4501000200089400007200D0020008000000144C4800000200BC228404020080",
INIT_15 => X"0010000104001000010440080000822900000000801010500A13404111008000",
INIT_16 => X"D1A0CA0000984D06403600086591900224002000400440104001040010000104",
INIT_17 => X"8DA368DA3685A1685A1685A1685A1685A1685A1685A1685A1685A1685A120D08",
INIT_18 => X"5A1685A1685A1685A1685A1685A368DA368DA368DA368DA368DA368DA368DA36",
INIT_19 => X"000000000000685A168DA368DA368DA368DA368DA368DA368DA368DA1685A168",
INIT_1A => X"6C20080AB9A28724904120E1999E91BCD151200802001038E2550A0010100000",
INIT_1B => X"68341A0D14514514514514514514514514514514514514534D34D34D34D344A1",
INIT_1C => X"268341A0D069349A0D069349A0D068341A4D268341A4D268341A0D068341A0D0",
INIT_1D => X"00000000000000000000000000000000000003FFFFFFFFFFFFFF8A6AC8341A4D",
INIT_1E => X"C2000557FEABEFA2D1400AA5D2AAAA00F7FFEAA10F7D17FFFFAAAE8000000000",
INIT_1F => X"03DFEFF7FFE8ABAF7802ABEFAAAE820000000021EFAA843DE00F7803FEBAFFFF",
INIT_20 => X"843DE00557BEAABAA2AEAABEFF78015555AA80174105555421EFF78028BEF5D0",
INIT_21 => X"504175FF0851401455555555EFA2FBC01FFF7AAAAB45557BC0155007FFDEBAAA",
INIT_22 => X"552A974AAA2843DEAA5D2A820BA000428AAAAA84154AAA2AA955FF00043DE005",
INIT_23 => X"AF7D1400BAAAAE821EFF7D17DEAA5D2AAAAAA5D557DE105D2EBDF55557FFDE00",
INIT_24 => X"BAFF803DF45FFD17DFFFFFD56AA00557FC201000517FFEFAAAEBDF45FFAEA8AB",
INIT_25 => X"FD7A2A48000000000000000000000000000000000000000000002ABFFA280154",
INIT_26 => X"AE38FF843DEBAEBFFC20285D75EFBC7A2DB400824120ADA38E3F1EFA28F7DF7D",
INIT_27 => X"421C7FF8028BEF41003FFD7F7F1EDA82F78E2DBD7A2A482038000A001C7A2803",
INIT_28 => X"1C716D1475FFEAAA28E3FE385D71E8AAAAAA0A8BC7EB8417555AA84104385D55",
INIT_29 => X"AA955C708003FE285D00155FF0055451555D5F575C7A2FBC51EFEBA0A8B6D557",
INIT_2A => X"12EBFF45497FFFE105D2E97482AA8038EAA412E850AA1C0428ABAB68E124BAA2",
INIT_2B => X"B6A0BFF55F7AEAAA82FFDF40092B6A4871EFFFD57FE825520ADA92495B7AE104",
INIT_2C => X"0000028BEFA28E124AAF7843AF7DEBDB78FFFE3DF6DA284175C001000557FFEF",
INIT_2D => X"AAA2D57FEAAF7FBFDF45AA800000000000000000000000000000000000000000",
INIT_2E => X"0BA082E82155AA802AAAAFF803DEBAAAFBC20BA55517DF55A2FBC201008003DE",
INIT_2F => X"5545A284000BA5D5340145F78028BFF08003DF45FFD57FE00FFAABFF45AA8002",
INIT_30 => X"D75FFA2842ABFF5555575FF55557FEAAA2AABFEAA5D5568ABAA2842AB55A2801",
INIT_31 => X"028ABAF7AA820BAAAAE9754500043DEBA5D04175EF0855575455D7BD5555A2FB",
INIT_32 => X"003DE00007FEAA10002ABFF450079FFE005D2A97400A2802AABA002A954AA5D0",
INIT_33 => X"0514200008517DFEFFF803FF45FFAAA8A00F7FBC2010FF80155EFF7D57DE005D",
INIT_34 => X"000000000000000000000028BFFA2AE820AAFF802ABEFAAFFEABEFAAFFFDEAA0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000200000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10044B00018248A2840112C00002C18000202300500030B3132000400992006",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110204",
INIT_02 => X"0801080200100000046558040080000041000000002402400800000009008010",
INIT_03 => X"00020201040000D0842242024210810802006400088000003080054288C10000",
INIT_04 => X"0000400088020000003020002000001002A0E881108032100002000800203040",
INIT_05 => X"04092A081000411841480001000000201000012800400010001081C040402000",
INIT_06 => X"10100001220001E0001802002020240208000369001520080100100909000266",
INIT_07 => X"4000220440020000090C0810210A040004A0410000C0000810000C4901036008",
INIT_08 => X"0000802100100140004200808809000C002000000000010F8102041320000000",
INIT_09 => X"2000000000000200828888800808000410800840100220211850004442004048",
INIT_0A => X"240A80800442400004C0010000060210200008B2022304880800410000200801",
INIT_0B => X"0000010008008020020100008000400120800004004821202001A05A00040180",
INIT_0C => X"08101400000000A01004101400000000A0100000081300410402080080003000",
INIT_0D => X"04101080000000A01004101080000000A0100540000040000000000000405100",
INIT_0E => X"00000040A80009000180000000000000004608004200040800000000000001A0",
INIT_0F => X"4000282000102000000080008000000000000000240800800140000040000000",
INIT_10 => X"00001A00000002000000000020013000100010080000000D0000040040000003",
INIT_11 => X"0000000021500000800010400000000000400900000088000000680000009000",
INIT_12 => X"008000800000000000086010000080000100000000000082C000100000200800",
INIT_13 => X"040004924040008020000200101100004000000000C019500050000800000000",
INIT_14 => X"4541008240801000804000108280800001001051A12481041080801010000080",
INIT_15 => X"4800048004480044800044000240022100884000901210440003C141102B088A",
INIT_16 => X"00044280009048485D4020080000140004046240020044000480044800448000",
INIT_17 => X"080200802008020080200802008020080200802008020080200802048026E011",
INIT_18 => X"0000000000000000000000000002008020080200802008020080200802008020",
INIT_19 => X"0000000000000080200000000000000000000000000000000000000000000000",
INIT_1A => X"CA83332A34488A8A28A29E195281FC1A72E24C2BF5A4D9555204428290100000",
INIT_1B => X"94CA65328A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A28A354",
INIT_1C => X"994CA6532995CAE572B94CA6532994CA6572B95CAE532994CA6532994CA65329",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF838CF1CAE532",
INIT_1E => X"7FFFFAAAE801FF08557DF4555516AA00007BEABEFAAD1555FFF7840000000000",
INIT_1F => X"56AA0000043FFEFA2FFFDE1008556ABEFA2D1400AA5D2AAAA00F7FFEAA10F7D1",
INIT_20 => X"84020000000021EFAA843DE00F7803FEBAFFFFC2000557FC0010AAD57FF45A2D",
INIT_21 => X"7FFE8ABAF7802ABEFAAAEA8BFF5D0415400F7FBFDEAA007FEAB45AAAE800AAF7",
INIT_22 => X"5D0415555557BFDFEF00517DE00A28028B450855421EFF78028BEF5D003DFEFF",
INIT_23 => X"A5D7FFDEBAF7AEBDE00557BEAABAA2AEAABEFF78015555AA80174105555401FF",
INIT_24 => X"FFF7AAAAB45557BC0155007FFDEBAAA8417410AAFFD7555AAD56AB45A2AE800A",
INIT_25 => X"5C7E380000000000000000000000000000000000000000000000155EFA2FBC01",
INIT_26 => X"DA38E3F1EFA28F7DF7DFD7A2A4801EF085F7AF6D55556AA381C75EABEFBED157",
INIT_27 => X"C0010AADF7AF6DB6D56FA3814003AFFFA2F1F8E381C516FBC7A2DB400824120A",
INIT_28 => X"5E8B45BEA0850BAE38002038000A001C7A2803AE38FF843DEBAEBFFC20285D75",
INIT_29 => X"8028BEF41003FFD7F7F1EDA82F78E2DBD7A2A4ADBEF550412428F7F5FDE92087",
INIT_2A => X"A84104385D55401C75504125455575FAFD7145578E10AA802FB450851421C7FF",
INIT_2B => X"BED56FB45BEA082082557BF8EBAF7AABFE385D71E8AAAAAA0A8BC7EB8417555A",
INIT_2C => X"00000175C7A2FBC51EFEBA0A8B6D5571C716D1475FFEAAA28E10438AAF5D2545",
INIT_2D => X"BA5D5568BEFF7D157555AA800000000000000000000000000000000000000000",
INIT_2E => X"F55A2FBC201008003DEAAA2D57FEAAF7FBFDF45AA80021FF007BE8BFF5D516AA",
INIT_2F => X"DEBAAAFBC20BA555140010AAFFE8BFFFFD17DEBA5D002ABFFA2D16AAAA55517D",
INIT_30 => X"020BAFFD17DE10005568B55FF80154BAA280020BA082E82155AA802AAAAFF803",
INIT_31 => X"43FF55085140145F78028BFF08003DF45FFD57FE00FFAABFF45AA803FFEF5500",
INIT_32 => X"842AB55A28015545A284000BA5D53421455504021555D556AB555D5568A00AA8",
INIT_33 => X"2AA800AAAAD142155F7D57DF45FF8002010557FEAAAAF7AABFEAA5D5568ABAA2",
INIT_34 => X"000000000000000000000015555A2FBD75FFA2842ABFF5555575FF55557FEAAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000023FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10180B05A0010402840602C2D001019000000300000000330A20080EC180002",
INIT_01 => X"AB400984B83008481800E0000C26426040000000080000088200000802112220",
INIT_02 => X"8801081438106400A4F55800008000004100000040CCE24208005000C9060032",
INIT_03 => X"00080D4912E6E440842254D002108153432004800880000030C0315688C00006",
INIT_04 => X"000048048002400048150000000002504230C899109032100020160880223000",
INIT_05 => X"040B2A229100410041088011100022201200012840440000B01088C0005C2400",
INIT_06 => X"287E4003225021C5021880C02000A40249048363A5992808110010090908022A",
INIT_07 => X"4044222987020C80152D8910210A0400252B74200045C86810000C5B0503286A",
INIT_08 => X"26509804400501400242C0B0B83B0134702000000000191FA162841324832069",
INIT_09 => X"3002000220001240820F8B2A08000040409018401001200159D80D64AA004041",
INIT_0A => X"020808852000420718C00101B0070310200008B60A23A51B2802467327200801",
INIT_0B => X"080802500C08832582810240812040912094068010050402214850444091019B",
INIT_0C => X"761B011986695014A96E1A8119865A5018C5A0A00012004104020808B0003000",
INIT_0D => X"AE1A811986695014A96E1B0119865A5018C5AF0062C38A4DB680A0D8241501D5",
INIT_0E => X"802CAB184E8F4101621B1BAC845542056A289A1BB2078A922DA2A8B180A2600A",
INIT_0F => X"392000224ACDE215883078681B5C05AA429189B60AC43CEC7F0272C3841DB528",
INIT_10 => X"51BCA1C90006C0C2958502861120C003104289A668B8CAB270106338317A3D94",
INIT_11 => X"A64090B89E015AAA880E48382EB8804B020A06020C67061BC785938085134CD5",
INIT_12 => X"C6284B2D20410AB4503089C00A8280819A5539D503336D61056ABA006282806C",
INIT_13 => X"060040142020015001004A00080042004000E8089C9003066E03513E41470126",
INIT_14 => X"4536708201C000908020349320008000A1000C09A9348498B000000000000080",
INIT_15 => X"32A0C32A0C32A0832A0C19504195040040000000801010028001400010010CBA",
INIT_16 => X"8104400000904C0C0964200841010954000444D280140050C32A0832A0C32A08",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090246811",
INIT_18 => X"1004010040100401004010040102409024090240902409024090240902409024",
INIT_19 => X"0000000000004010040100401004010040100401004010040100401004010040",
INIT_1A => X"488292A831308E0000000A11100830181621409A14E871104201400284000000",
INIT_1B => X"0000000000000000000000000000000000000000000000020820820820820A05",
INIT_1C => X"0000000402000000000000000000010080000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8C0F00000000",
INIT_1E => X"555FFF784020AAF7D542155F7D1400AAF7FFFDE00F7842AA00002A8000000000",
INIT_1F => X"A800AA007FFDFFFA28428A000000001FF08557DF4555516AA00007BEABEFAAD1",
INIT_20 => X"FBEABEFA2D1400AA5D2AAAA00F7FFEAA10F7D17FFFFAAAEA8ABAFFD17FEBAFFA",
INIT_21 => X"0043FFEFA2FFFDE1008556AB45555568A10A2FFC00AAF78028AAAFF84020AAFF",
INIT_22 => X"FFD1555FF0804000AA000428A10AAAA801EFFFD140010AAD57FF45A2D56AA000",
INIT_23 => X"FA2FBFFF550000020000000021EFAA843DE00F7803FEBAFFFFC2000557FC0155",
INIT_24 => X"00F7FBFDEAA007FEAB45AAAE800AAF78428B45A28428A10087FD7400552EBDFE",
INIT_25 => X"A101C2A80000000000000000000000000000000000000000000028BFF5D04154",
INIT_26 => X"AA381C75EABEFBED1575C7E380000BAF7DB4016DE3DF450AAF7F1FDE38FF8A2D",
INIT_27 => X"AFABAFFDF7AE82F7AA870AA0071F8FFFBE842DA101C0E001EF085F7AF6D55556",
INIT_28 => X"42DAAAE38A02082E3FBEFBC7A2DB400824120ADA38E3F1EFA28F7DF7DFD7A2A4",
INIT_29 => X"DF7AF6DB6D56FA3814003AFFFA2F1F8E381C516DB455D5B68A28A2FFC20AAEB8",
INIT_2A => X"BFFC20285D75C2145F7DF525EF140A050AA1C0028A28AAA4801FFE3DF40010AA",
INIT_2B => X"007FD74284120BFFFFBEF1F8F7D080A02038000A001C7A2803AE38FF843DEBAE",
INIT_2C => X"000002DBEF550412428F7F5FDE920875E8B45BEA0850BAE3802DB6DAA8A28A00",
INIT_2D => X"AAF7D57DEAAF7AABDE10552E8000000000000000000000000000000000000000",
INIT_2E => X"1FF007BE8BFF5D516AABA5D5568BEFF7D157555AA80020BAFFFBC01EFA2FFD74",
INIT_2F => X"FEAAF7FBFDF45AA803FEBAFFFBEAA00F7AE974BA085568BEFF7803FE10552E82",
INIT_30 => X"EAAAAA2FFC00AAAA803FEAAA2AA82000A2FFFDF55A2FBC201008003DEAAA2D57",
INIT_31 => X"0001FFAAFFC0010AAFFE8BFFFFD17DEBA5D002ABFFA2D16AAAA55517DF55557F",
INIT_32 => X"802AAAAFF803DEBAAAFBC20BA555142155F7FFC01EF552E974BA550028ABAA28",
INIT_33 => X"2803FFFFA2AAAAA00007FD74BA08003DFFFFFD16ABFF082E820BA082E82155AA",
INIT_34 => X"00000000000000000000003FFEF5500020BAFFD17DE10005568B55FF80154BAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000200000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A50080B01BC002006940202C0DE041196A83183000000023322287E0FC000006",
INIT_01 => X"0E000C068000E04D40238000001702684000000008000008820009280A553231",
INIT_02 => X"2809AD0E7D180040945008040090000061800000C0E2F66009DA3D11CB148015",
INIT_03 => X"421A0A0012F6F8D2108216E24842005B8A20640008800000B8E0141C28851006",
INIT_04 => X"02004000890200001837830011998C31C09060DC104000102002140900003548",
INIT_05 => X"0402002BC200009841090001200006200800000020480010A4100100001C2000",
INIT_06 => X"287FC003230001D0001806C0060CB0622000037085C820000000100C0C200008",
INIT_07 => X"CE64B663DFA314C803292140890C0601F472D1640051F80C10020C493F033432",
INIT_08 => X"67C081000111814004C20481A92940EA7A3020480000071F846890162E135038",
INIT_09 => X"240048108488024082488BAF08000020800629441004300421800F04F8000001",
INIT_0A => X"A0200E0BF40063FF9DC0010000180018200408B27E234913E900067F04D40C01",
INIT_0B => X"002002801000A04200000000000000000000029D204B7C0382FD0100F3F9F80F",
INIT_0C => X"7E0B348EDAC3900F6EFA0B158EDA93900F6EE230381208008001007A80001100",
INIT_0D => X"CA0B158EDAC3900F6EFA0B348EDA93900F6EE8421392C96B1237E0D8BD9628F9",
INIT_0E => X"412EDD2B47CFF812A383430C669E622DBC31D73F6006A5891533EF9500EAE64B",
INIT_0F => X"BA30E022DAD8C100CA39E8CEBE66C2B083798D341B10DE7E14400392C74CAEAD",
INIT_10 => X"71A9C5DD00B12728D5360234D62A49FAB442994B3238D4E2FB104636652E19B8",
INIT_11 => X"C800DA550C29F36A8A2554E48A6430469392526208C6CC95C33717D885329664",
INIT_12 => X"51B60585A5C28895962502E9F36A828C4999AF580395542D27CDBA0020F0FABA",
INIT_13 => X"0000001E404011F066000A000EE040000000873FB80B8A00EF03F56CC12B416A",
INIT_14 => X"4D667C06CC6816B300403C13E2000000460010400000010CE080801010000080",
INIT_15 => X"72F0C72F0872F0872F0C597863978421040800209010124ACA03414158228430",
INIT_16 => X"00104280A89A4D004000000800001D5E05182493C5BC5AF0872F0C72F0872F08",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000010000",
INIT_18 => X"8020080200802008020080200800000000000000000000000000000000000000",
INIT_19 => X"0000000000000080200802008020080200802008020080200802008020080200",
INIT_1A => X"E02000028DCA05A8A28A2048C1111026C152A2316246000CB054420210100000",
INIT_1B => X"C864321904104104104104104104104104104104104104124924924924924481",
INIT_1C => X"2C964B2592C964B2592C964B2592C964B2592C964B2592C964B2190C86432190",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800FFD64B259",
INIT_1E => X"2AA00002AAAA10FF8002155F7FFC2000080417555FFAA80155F7840000000000",
INIT_1F => X"FE8AAA080000155F7FFFDEAA0000020AAF7D542155F7D1400AAF7FFFDE00F784",
INIT_20 => X"2E801FF08557DF4555516AA00007BEABEFAAD1555FFF7842AB55080000145557",
INIT_21 => X"07FFDFFFA28428A00000028B4555043DFFFFFAE82000FF80020AAA2AAAABFF00",
INIT_22 => X"A284174AAFF8428AAAFF8415545AAFBD7545F7AAA8ABAFFD17FEBAFFAA800AA0",
INIT_23 => X"5F7FFFDEAA08556ABEFA2D1400AA5D2AAAA00F7FFEAA10F7D17FFFFAAAE80000",
INIT_24 => X"10A2FFC00AAF78028AAAFF84020AAFFFBC21550800000105D55400AA082A8215",
INIT_25 => X"145F7840000000000000000000000000000000000000000000002AB45555568A",
INIT_26 => X"50AAF7F1FDE38FF8A2DA101C2AAFA00EB8E0516DE3F5C000014041256DEBA487",
INIT_27 => X"2FB551C0E0516D417FEDA921C000017DEBF5FDE92080E000BAF7DB4016DE3DF4",
INIT_28 => X"0070BAAAAAADBD70820801EF085F7AF6D55556AA381C75EABEFBED1575C7E380",
INIT_29 => X"DF7AE82F7AA870AA0071F8FFFBE842DA101C0E2DB55410A3FFC7F7A087000FF8",
INIT_2A => X"7DF7DFD7A2A480000BE8A17482F78A28A92E3841556DA2FBD7545F7AAAFABAFF",
INIT_2B => X"41554508208208017DF7F5FDE9208556FBC7A2DB400824120ADA38E3F1EFA28F",
INIT_2C => X"000002DB455D5B68A28A2FFC20AAEB842DAAAE38A02082E3FBC217D1C0E05000",
INIT_2D => X"005504001FFAA8015545F7800000000000000000000000000000000000000000",
INIT_2E => X"0BAFFFBC01EFA2FFD74AAF7D57DEAAF7AABDE10552EBDE00AAAE975FFAAD1420",
INIT_2F => X"8BEFF7D157555AA803DF45552E975EF007FFFE005504001FFAAD17DE00082E82",
INIT_30 => X"BFF55FF8017410FF84154BAAAAABFF450000021FF007BE8BFF5D516AABA5D556",
INIT_31 => X"BD5555F7AEBFEBAFFFBEAA00F7AE974BA085568BEFF7803FE10552EBDF45002E",
INIT_32 => X"003DEAAA2D57FEAAF7FBFDF45AA8002000FFAE95400F7AEA8A10A284175FFAAF",
INIT_33 => X"2FFC21EF552A954100851554000004021FFFFD17DE1008517DF55A2FBC201008",
INIT_34 => X"00000000000000000000003DF55557FEAAAAA2FFC00AAAA803FEAAA2AA82000A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10110A0441812402840402822007818000E00700000000330A3000000008042",
INIT_01 => X"A1400984B830C848180260000C0042404001000008220008A200100802110200",
INIT_02 => X"88010C02801040002475580400800000410000000064024608134C0CC9018034",
INIT_03 => X"00020201926220D084234212421085084300648A0880000630C0654288C10000",
INIT_04 => X"00104884880A4400403000004800027102A0E88110D83210642EA809C0203040",
INIT_05 => X"04092A08138041184109C001380000201A008128044E00754010C9C192D82400",
INIT_06 => X"201800012372A1D72A180000204024024954A3670819290951001009092C0222",
INIT_07 => X"4000220B40020C80052C0A12292A040005715540015E006810001C4B01032C7E",
INIT_08 => X"9032881000140140024200808839005C002010800000155F8122851320016400",
INIT_09 => X"2C80080200801280825A988008000040008208401005B3071859006442004054",
INIT_0A => X"200810940400720005C0030192072310200028B6022346080802E001A5600801",
INIT_0B => X"206822F20CA8826AC2A14250A128509528954404144C200425010040000001B0",
INIT_0C => X"A41AA5B7344C10B383081BA4B7341C10B3831034081200000000000430003000",
INIT_0D => X"381BA4B7344C10B383081AA5B7341C10B383110218CB0E54C2EA404A4F03D404",
INIT_0E => X"A008E730A01AB113A5524E6ACA678001CE3E20A5B284ED1132909C72885A2B2C",
INIT_0F => X"6430202021252991C22C99731014AC3CC0C0B8182597A801610218CB0C3548B3",
INIT_10 => X"5194332B018A444AEA2701288A15A151EC5952E44128CA194517354C180A3C06",
INIT_11 => X"D50048A411C158BB0A7910142C771804C8A0ADA2E6A983014780CA28B2A5C882",
INIT_12 => X"F8BE8E3E1E0109472C3EB50158BB02D09852745F80112C428562EE0353635232",
INIT_13 => X"02414032646000826080C20001104240480068001C9B9150A0000297046E4023",
INIT_14 => X"4510008241C80290882400908000A000A1000809A93485D61000000000000080",
INIT_15 => X"00000000040000000000000020000000000000008010102A82014100101118BA",
INIT_16 => X"A10441010090480C096420184321040002844840000000004000000000400000",
INIT_17 => X"0942509425094250942509425094250942509425094250942509425094246A10",
INIT_18 => X"9425094250942509425094250942509425094250942509425094250942509425",
INIT_19 => X"0000000000005094250942509425094250942509425094250942509425094250",
INIT_1A => X"BFBFBFBF7DDF3BAAAAAABEFDDFE7EFBEFFE7CFC3F7EFFF7DF7E24502A8000000",
INIT_1B => X"F5FAFD7EBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAFFD",
INIT_1C => X"BF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EB",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800FFDFAFD7E",
INIT_1E => X"80155F7842AB55552E821FFFFD5555EF552ABDFEF007FE8A00AAFBC000000000",
INIT_1F => X"BD55EFAAD1554BA00556AA00AAD16AA10FF8002155F7FFC2000080417555FFAA",
INIT_20 => X"55420AAF7D542155F7D1400AAF7FFFDE00F7842AA00002A821EF5D7BC21FFFFF",
INIT_21 => X"80000155F7FFFDEAA00002AB45082A821EF5D557FF45A2AABFEBA082A975555D",
INIT_22 => X"A2FFE8BEF5D517FF455D554214500043DEBAAAFFEAB55080000145557FE8AAA0",
INIT_23 => X"0552EBFEAAAAD1401FF08557DF4555516AA00007BEABEFAAD1555FFF7842AABA",
INIT_24 => X"FFFFAE82000FF80020AAA2AAAABFF002E80000AAAABDF555D2E955EFA28428A1",
INIT_25 => X"A28AAF5C0000000000000000000000000000000000000000000028B4555043DF",
INIT_26 => X"000014041256DEBA487145F78428B6D4120851FFEBD5525C74124B8FC71C71EF",
INIT_27 => X"871C74975C01FFEBF5D25EFA2D555482085F6FA28AAD16FA00EB8E0516DE3F5C",
INIT_28 => X"0BFE921C2E9557D415B400BAF7DB4016DE3DF450AAF7F1FDE38FF8A2DA101C2A",
INIT_29 => X"0E0516D417FEDA921C000017DEBF5FDE92080E2AB7D1C24851FF495F7FF55A2A",
INIT_2A => X"ED1575C7E38028A82B6F1E8BFF495F78F7D49554214508003FEAABEFFEFB551C",
INIT_2B => X"5D20905C7AA842DA00492EBFEAABED1401EF085F7AF6D55556AA381C75EABEFB",
INIT_2C => X"000002DB55410A3FFC7F7A087000FF80070BAAAAAADBD7082087000AAA4BFF7D",
INIT_2D => X"4508042AB455D517DEBAA2D54000000000000000000000000000000000000000",
INIT_2E => X"E00AAAE975FFAAD1420005504001FFAA8015545F78028BFF0004175EFA2D5421",
INIT_2F => X"DEAAF7AABDE10552E975450051401EFA2D5421EFAAD557410007BFDEAAA2D57D",
INIT_30 => X"175FF087BFFF45AA843FE005D2A955FF087BC20BAFFFBC01EFA2FFD74AAF7D57",
INIT_31 => X"03FEBAFFFBFDF45552E975EF007FFFE005504001FFAAD17DE00082EA8BFF5504",
INIT_32 => X"516AABA5D5568BEFF7D157555AA8028A00FFD16ABFF087BEABEF005542155000",
INIT_33 => X"00017410AA803DFEF550402155A2843FE00082ABFEAAFFD5421FF007BE8BFF5D",
INIT_34 => X"00000000000000000000003DF45002EBFF55FF8017410FF84154BAAAAABFF450",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000033FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10020A000180000284008280000281800000030000000033022000000580002",
INIT_01 => X"A140098018300848184860000C20C24040000000084000084200000000110200",
INIT_02 => X"88010C5A8010A600A4F558040080000041000000022C024008003CCCC9028030",
INIT_03 => X"0002074F200904D0842242024210810803006480088000003081054288C10000",
INIT_04 => X"0000480488024000403000000000001002A0E881108032100002000800203040",
INIT_05 => X"04092A081000411841080001000000201000012800400010001081C000402000",
INIT_06 => X"80500001221021C1021800002000240249048361001128081100100909000222",
INIT_07 => X"4000220050020480152D0A142D0A8400043B45400040006810000C5901033D78",
INIT_08 => X"0010880000100140024280808829029C002000000000053FA142051324902030",
INIT_09 => X"2000000000000200820888800800004000800840100020011858006442004040",
INIT_0A => X"200800840400400005C0010190070310200008B202236D080802400001600801",
INIT_0B => X"000000100C088020028102408120409120940404104C20002101004000000110",
INIT_0C => X"5210040000B0E0A0000210040000E0E0A0000190081200000000000000003000",
INIT_0D => X"0210008000B0E0A0000210008000E0E0A0000B02740421A0E5D1A02400205080",
INIT_0E => X"40110080A4006110510C14D18178E01200860008920106460D4501CB00011130",
INIT_0F => X"411420220080220C0093C38923240ABBC00905C33C6000400F02740412C0715C",
INIT_10 => X"8000120800658992F3C700C3018120000041DB011CC000090012565306500002",
INIT_11 => X"E240240A8340000200067EAA8CB65809240C09024A4AE0CA0000480083968239",
INIT_12 => X"7DB0D0200900422ACA4B28000002002B46867DBC002A830280000800F7B7A0B1",
INIT_13 => X"020040126060008020000200000042004005800004801150A00341244000845C",
INIT_14 => X"4500008240800000802000908000800001000009A92481041000000000000080",
INIT_15 => X"000040000000000000040000000000000000000080101000000141001001088A",
INIT_16 => X"810440000090480C096420084101040000044040000000004000040000000000",
INIT_17 => X"0902409024090240902409024090240902409024090240902409024090246810",
INIT_18 => X"9024090240902409024090240902409024090240902409024090240902409024",
INIT_19 => X"0000000000004090240902409024090240902409024090240902409024090240",
INIT_1A => X"EFBBBBAABCDABF9E79E7BEF9CB91FE1EF7D3AEB9F3E6FF7DF650400280000000",
INIT_1B => X"FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E7FC",
INIT_1C => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8FF000FE7F3F",
INIT_1E => X"E8A00AAFBE8BEFA2D568ABA00003DF555555574AAAAAEAAB45082E8000000000",
INIT_1F => X"02AABA555155400557BC2010557BEAB55552E821FFFFD5555EF552ABDFEF007F",
INIT_20 => X"002AA10FF8002155F7FFC2000080417555FFAA80155F78428AAA007FE8A10080",
INIT_21 => X"AD1554BA00556AA00AAD140145AA8028ABA002EBFFFF082EBDEBAA2D1420105D",
INIT_22 => X"A2AEA8A10080428A10FFAEBFFEF5D0428B45A2FFC21EF5D7BC21FFFFFBD55EFA",
INIT_23 => X"5F7FBC0010FFAA820AAF7D542155F7D1400AAF7FFFDE00F7842AA00002A80155",
INIT_24 => X"EF5D557FF45A2AABFEBA082A975555D55400BA005568A000000175FFF7D15554",
INIT_25 => X"B6D00248000000000000000000000000000000000000000000002AB45082A821",
INIT_26 => X"25C74124B8FC71C71EFA28AAF5E8BFFB6D56DA82000E38F6D4155504AAA2AEAA",
INIT_27 => X"28ABA147FEDA10080E2AAAA555552400417FC20005D75E8B6D4120851FFEBD55",
INIT_28 => X"4BAEAAB6DB4202849042FA00EB8E0516DE3F5C000014041256DEBA487145F784",
INIT_29 => X"75C01FFEBF5D25EFA2D555482085F6FA28AAD147155BE8028A82002EB8FC7002",
INIT_2A => X"F8A2DA101C2A80145B6AEA8A10080E2DA00F7A0BDFD7550428B55A2F1C71C749",
INIT_2B => X"0004175FFE3D15757DE3F5C0038FFAA800BAF7DB4016DE3DF450AAF7F1FDE38F",
INIT_2C => X"000002AB7D1C24851FF495F7FF55A2A0BFE921C2E9557D415B400AA00556DA00",
INIT_2D => X"EF0051400AAA2AAAABFF08000000000000000000000000000000000000000000",
INIT_2E => X"BFF0004175EFA2D54214508042AB455D517DEBAA2D568BEFFFD57FE10002AAAB",
INIT_2F => X"01FFAA8015545F78028AAA557FFFE00082EAAAAA5D5142000007BC20105D5568",
INIT_30 => X"28A00082EAAB45000028ABAFFFBC20AA08043DE00AAAE975FFAAD14200055040",
INIT_31 => X"02AB55AAD1575450051401EFA2D5421EFAAD557410007BFDEAAA2D557555FF80",
INIT_32 => X"FFD74AAF7D57DEAAF7AABDE10552E82155FFAAA8A10002ABFE00F7803FF555D0",
INIT_33 => X"87BC20AA00517DE000804175EFAAD1555EFA2D1420BAFFAE820BAFFFBC01EFA2",
INIT_34 => X"000000000000000000000028BFF5504175FF087BFFF45AA843FE005D2A955FF0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A10000A000000000284000280000001800020030000000033022000000180002",
INIT_01 => X"A140098018300848180060000C00424040000000080000080200000000110200",
INIT_02 => X"080108000010E60004E55800008000004100000000040240080000C009170016",
INIT_03 => X"0000000100000040842240000210810002000400888000003080014288C00000",
INIT_04 => X"000440009282000001100000000000100220C8811080321000000228002A3000",
INIT_05 => X"04092A0010004300418800510000A6201000012A64400000145080C000422000",
INIT_06 => X"00100001220001C00018821020402402080003772019200001001009090002AA",
INIT_07 => X"4000220000021840010C8912250A0400042044400040006810000C4901032B18",
INIT_08 => X"0022810000058140024280A0A8190004002030C00000016F8122041320000000",
INIT_09 => X"20000000000002C0820888008800000000800840100020011850004402004040",
INIT_0A => X"00080094000062000180010180060210200008B2022304080800400003E00801",
INIT_0B => X"0000000008008020020000000000000100800000000000002500004000000130",
INIT_0C => X"0010108000000000000010108000000000000230001200000000000420003000",
INIT_0D => X"0010140000000000000010140000000000000100000040000000000000000000",
INIT_0E => X"0000000000000100008040000000000000000000020000090000000000000000",
INIT_0F => X"0030002000406000000000068409014000000000000000000100000040000000",
INIT_10 => X"0000000800000201000800000000000000400048000000000010000440000000",
INIT_11 => X"00A0000000000002000000441108800000000002008008000000000080201000",
INIT_12 => X"0242038B82800000000000000002000001000000000000000000080000001844",
INIT_13 => X"000000100000000005C04A000000400000000000000001062000000400000000",
INIT_14 => X"4500008200800000800000100000800001000001A12480001000000000000080",
INIT_15 => X"000000000000000000040000200002000000000080101000004140001001088A",
INIT_16 => X"0004400000904808094020080000000000044040000000004000040000400004",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000046000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000400280000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000000000",
INIT_1E => X"AAB45082EBFE000004020AA552E80000F7FBC214555003DE10A2FBC000000000",
INIT_1F => X"BE8A10F7802AA0055003FE10007BE8BEFA2D568ABA00003DF555555574AAAAAE",
INIT_20 => X"AEAAB55552E821FFFFD5555EF552ABDFEF007FE8A00AAFBFDEBA555568BEFA2F",
INIT_21 => X"55155400557BC2010557BFFFEFA2FFC20005D2A955EFF78428BEFAAD17DF55AA",
INIT_22 => X"5D2AA8B45AAD57FF55A2FBC21FFA28415400FF8028AAA007FE8A1008002AABA5",
INIT_23 => X"A002E9740055516AA10FF8002155F7FFC2000080417555FFAA80155F7843DF45",
INIT_24 => X"BA002EBFFFF082EBDEBAA2D1420105D003FFFF08514200055002AA00AA802AAB",
INIT_25 => X"E28B6FFC0000000000000000000000000000000000000000000000145AA8028A",
INIT_26 => X"8F6D4155504AAA2AEAAB6D0024B8E381C0A00092412A87010E3F5C0145410E3D",
INIT_27 => X"F8EAA495F68BFFA2F1EFA38E38428A005D0038E28147FE8BFFB6D56DA82000E3",
INIT_28 => X"428BEFB6DB7DF45AAAEA8B6D4120851FFEBD5525C74124B8FC71C71EFA28AAF5",
INIT_29 => X"7FEDA10080E2AAAA555552400417FC20005D75F8FFFBEF5C0000492A955FFF78",
INIT_2A => X"BA487145F7843FF7D4120A8B6DAAD17FF55B6F5C21EFAA8E10400E38E28ABA14",
INIT_2B => X"41002FA38A2842AA82142095428415F6FA00EB8E0516DE3F5C000014041256DE",
INIT_2C => X"0000007155BE8028A82002EB8FC70024BAEAAB6DB4202849043FFC7005F45010",
INIT_2D => X"00A2D542155002ABDEBAF7FBC000000000000000000000000000000000000000",
INIT_2E => X"BEFFFD57FE10002AAABEF0051400AAA2AAAABFF08002AAAA5D2A82000082E954",
INIT_2F => X"AB455D517DEBAA2D56AABA087BEABEFAAD57DEAAA2802AA105D002AABA5D7BE8",
INIT_30 => X"42010082A955EFFF8428BFFFFFBFDF55A2AEA8BFF0004175EFA2D54214508042",
INIT_31 => X"A82000AAAAA8AAA557FFFE00082EAAAAA5D5142000007BC20105D556ABFFF7D1",
INIT_32 => X"D1420005504001FFAA8015545F7803FFEF08002ABEFA2D57DF45F7D1401FFA2A",
INIT_33 => X"8043FF55087BD740000043DEAAA2842AA005D00154AA007BFDE00AAAE975FFAA",
INIT_34 => X"000000000000000000000017555FF8028A00082EAAB45000028ABAFFFBC20AA0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000300000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA22C618B1000482B688B186588884862A400438255FC38381441205BA803003",
INIT_01 => X"8645A80028404C211203A952A90341080B173340412000E1005D628000820484",
INIT_02 => X"A101A9006DC1084833011850AAC55001349B10881802821808B4110007005E11",
INIT_03 => X"0202115002BB10080080006020020001A61036202800000D2410104200404550",
INIT_04 => X"2FE962000017102918900948514522CE09200C0D590569398ADBF8CC1E50E480",
INIT_05 => X"5E6023002834854AE41C1E8782F508F2A15B71D412E0AFD9C2990DA56FF0B55A",
INIT_06 => X"B9B9E55402000340003200220A86012D0000000480D0400001555960540180A0",
INIT_07 => X"40D890101DBD400901442800817C2901F400868554DE240000A80090CE82A803",
INIT_08 => X"0122004000005665510320C9C90510025A8A00000A0A048F550A440E0001380C",
INIT_09 => X"2060410280081116C8204D016CB2CB290008008279580411289000000118A905",
INIT_0A => X"00008176802203180025699200140001A15000017F0051D0F837324E002A8A56",
INIT_0B => X"4485D000000124002400000000000001004010A8812831605DA0000A054052E4",
INIT_0C => X"B5320018CAC99BA0A3B9320018CAAAADA0C343F1AC1B01040A00202489551455",
INIT_0D => X"59320018CAC99BA0ACB9320018CAAAADA0CC421CA003B694B68018FAAA708E2C",
INIT_0E => X"B2449A3FF2FA04E5E09B128834ADB1443A1891E4A928C29020E6A8524CE7A3EE",
INIT_0F => X"2375B801324301AB0067622E5E5404B2A5A40B1E6644AF0F021EA003AC24352A",
INIT_10 => X"0A8C241815FEB6A9158863F638FB60ED838E890B703C6260D8E3A21275714C90",
INIT_11 => X"15F11133D171727A2550EE2F1BA0064F70DBDB1C74424E91E1C194C71D1216F5",
INIT_12 => X"432A2B2D001F803471A9A960E57245FDF9D364DBD9435A6D45C9E81BED555E4C",
INIT_13 => X"C00006B0800000038814B72AB01508150013F162119014204373517700ACCC59",
INIT_14 => X"300208092B940192D1000000000000A8A5AA80018120E00066000000000012CA",
INIT_15 => X"1000110001100011000108000880008000520228080108039501200848002912",
INIT_16 => X"081500008A422150884081AC9000010003561180063DB4F61100011000110001",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000012000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"BCBF0F2C688A8D3CF3CF0A7A898D21B4C9838D3030EF5168A360400000000000",
INIT_1B => X"E9F47A7D345345345345345345345345345345345345345145145145145147A5",
INIT_1C => X"3E9F4FA3D1E8F47A3D1E8F47A3D1E9F4FA7D3E9F4FA7D3E9F4FA7D1E9F47A7D1",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800001F4FA7D",
INIT_1E => X"3DE10A2FBC21FFFFFBFDF45A2D56AB45FFFFD54BAFF80001FF002A8000000000",
INIT_1F => X"FFFE005D7BC0010002E954AA087FFFE000004020AA552E80000F7FBC21455500",
INIT_20 => X"FFE8BEFA2D568ABA00003DF555555574AAAAAEAAB45082E974BA5D7BFDF55A2F",
INIT_21 => X"7802AA0055003FE10007BC0000082A97400550017410FFD1555550000020BAAA",
INIT_22 => X"AAFBD74105504021FF5D2EAAABAFFFBD55FF002ABDEBA555568BEFA2FBE8A10F",
INIT_23 => X"0007FC00AA087FEAB55552E821FFFFD5555EF552ABDFEF007FE8A00AAFBD55EF",
INIT_24 => X"005D2A955EFF78428BEFAAD17DF55AAAE820AA5D517DF45AAFFFFEAAFFAABFE1",
INIT_25 => X"1FF08248000000000000000000000000000000000000000000003FFEFA2FFC20",
INIT_26 => X"7010E3F5C0145410E3DE28B6FFC21C7E3F1F8F55AADB6FB6DFFFBD54AAE38E02",
INIT_27 => X"92482497BFDF45AAFFF8E385D7BC5000002E904BA1C7FF8E381C0A00092412A8",
INIT_28 => X"B555450804070BABEF5E8BFFB6D56DA82000E38F6D4155504AAA2AEAAB6D0024",
INIT_29 => X"5F68BFFA2F1EFA38E38428A005D0038E28147FC2010142E90428490015400FFD",
INIT_2A => X"C71EFA28AAF5D25D7B6F1D54384904021FF5D2AADAAAFFF1D55FF002EB8EAA49",
INIT_2B => X"A2F1FDEAAEBAABDE001471C20921475E8B6D4120851FFEBD5525C74124B8FC71",
INIT_2C => X"0000038FFFBEF5C0000492A955FFF78428BEFB6DB7DF45AAAE820925D5B7DF45",
INIT_2D => X"EFF7FFD54AAAAAA801EF00000000000000000000000000000000000000000000",
INIT_2E => X"AAA5D2A82000082E95400A2D542155002ABDEBAF7FBC2145AAD568B45AAFBFFF",
INIT_2F => X"00AAA2AAAABFF080000000087BFDF55A2FFE8AAA557FD7410082A800AA557BEA",
INIT_30 => X"800BA080417400F7FBD75450800174AAFFD168BEFFFD57FE10002AAABEF00514",
INIT_31 => X"1575EF082EAAABA087BEABEFAAD57DEAAA2802AA105D002AABA5D7BC20005D2E",
INIT_32 => X"D54214508042AB455D517DEBAA2D540155F7D1554AA0800001EF5D2ABDEBAF7D",
INIT_33 => X"2AE82010557FFDF55A2D57FEAAAAAEBFE10555140000555568BFF0004175EFA2",
INIT_34 => X"00000000000000000000002ABFFF7D142010082A955EFFF8428BFFFFFBFDF55A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000100000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5284CE4FB7BD2C8994A13392DBD02E14006B82AC7E800D44D3DD2FD5F9B961C0",
INIT_01 => X"F8ACD01F7E03FC6793F2199B39FC233C11D93AE6F3BB92B32091DBC339B24542",
INIT_02 => X"8F333007FD6808092A2AFA6667033DB50853379C10BFF70F1BD011110F205F18",
INIT_03 => X"5295B6957FCBE0DAD63ABF836B58EAFE060478202022234B2E0303FDC9E18339",
INIT_04 => X"6DE90201BF90102103AF158E805428249851BFB2C106592088DBF8400A5055C2",
INIT_05 => X"3824BD7F80148D9E07100A8201ED01C1A19B68F40A807ED9C18114956FF081DB",
INIT_06 => X"6A8F033DD800000000050716BE9F57F8AC000807DFD9B00000CF20E5E1818B1B",
INIT_07 => X"86481240FE05A109228E2C0891D772A6F40045B8CF30E085DD2ED57D4EED08CA",
INIT_08 => X"DF23800005981C0338190549C904182B6113870022000488C08B46268A001508",
INIT_09 => X"823DF78CDB6CA60E0E28EFFE2061872F80C1684A80C8604085F0074D3B72637F",
INIT_0A => X"BD2FAD7FE653C3BA1FF33E0E001E000B3A5DAADAFDDA5DA79350CFB8013E7437",
INIT_0B => X"C5C3D00018006C681700000000000000020012E9E10A31EB5FF9296A67F5B4FF",
INIT_0C => X"542A6FEEB2533EA160782A6FEEB2333EA16031F2BD47BDA2CA5D8164FCCFE833",
INIT_0D => X"F82A6FEEB2533EA160782A6FEEB2333EA160391BEFF2C32FB695F919110D5ECE",
INIT_0E => X"5A86840354D1706FFFA3EF6E24B6D18C0D06638A207CFDE1F7DDAD76D5282400",
INIT_0F => X"4D77FAAB77CE3AF3EE78F58DB737E6E43E59AFE4A59B57679D19EFF2C7573FAD",
INIT_10 => X"72CA52606DFED6CA55334C04C04FF7D7A0ABD6DAAAB96529382B74E4E1FE4ACA",
INIT_11 => X"AA1A184045D5D7A870D2F5A5D7522D1281017F056E9C9C3FC95949C157ADB555",
INIT_12 => X"A58949D5B5C85F97871876F7D7E859FDEB974F486905001FDF5FA0D719F9956E",
INIT_13 => X"70021EE341036BF368128419FB5560158015177F916A039EF41FDB34A91F432E",
INIT_14 => X"1D0A7CC9AE7A08BFF0001D35682AC0CE8FCCC200A59BDD2FFE3F3EC7C7DEF206",
INIT_15 => X"BCF4FBCF4FBCF4FBCF4FBE7A7DE7A7800617112E46F05D02DD814102F800633F",
INIT_16 => X"00179C16DECF67F08BC02F9086000D9E8A3F06ABD73DBCF4FBCF4FBCF4FBCF4F",
INIT_17 => X"000000000000000000000000000000000000000000000000000000000005F080",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"930D0D1B9000303AEBAE88BE013DB9880A5D25C0408006114F981800C0000000",
INIT_1B => X"351A8D069A6BAE9A69A6BAE9A6BAE9A69A6BAE9A6BAE9A69A69A69A69A69A918",
INIT_1C => X"A351A8D46A351A8D46A351A8D46A341A0D068341A0D068341A0D068351A8D068",
INIT_1D => X"00000000000000000000000000000000000003FFFFFFFFFFFFFF8000011A8D46",
INIT_1E => X"001FF002A821FFFFFFFFFFFFFFBFDFEFAAD142010007BEAB55FFAA8000000000",
INIT_1F => X"A975EFA2D140145007BC21FF5D2A821FFFFFBFDF45A2D56AB45FFFFD54BAFF80",
INIT_20 => X"7BFFE000004020AA552E80000F7FBC214555003DE10A2FBEAB45A28000010082",
INIT_21 => X"D7BC0010002E954AA087FD7400082E954AA0800154AA0855575FFAAD57FE005D",
INIT_22 => X"F7D16AB45FFFFEABEF007BD74005555555EFF7AE974BA5D7BFDF55A2FFFFE005",
INIT_23 => X"5555568B45552EA8BEFA2D568ABA00003DF555555574AAAAAEAAB45082EBFFFF",
INIT_24 => X"00550017410FFD1555550000020BAAAFFC0145AA84154BA082E801FFAAFBC015",
INIT_25 => X"B7DEBA480000000000000000000000000000000000000000000000000082A974",
INIT_26 => X"FB6DFFFBD54AAE38E021FF0824851FFFFFFFFFEFF7F1FAFD7A2D5400001C7BED",
INIT_27 => X"EFB45AA8E070281C20925FFBEDB451451C7BC01EF4124821C7E3F1F8F55AADB6",
INIT_28 => X"5505EFBEDB7AE385D7FF8E381C0A00092412A87010E3F5C0145410E3DE28B6FF",
INIT_29 => X"7BFDF45AAFFF8E385D7BC5000002E904BA1C7FD54280024924AA1404174AA005",
INIT_2A => X"2AEAAB6D0024BFFD7FFDB6AB7DFFF5EDBC71C7BD54005D5B575EFEBAE9248249",
INIT_2B => X"1C20801FFB6F5C0145555B68B7D4124A8BFFB6D56DA82000E38F6D4155504AAA",
INIT_2C => X"0000002010142E90428490015400FFDB555450804070BABEF5C516DAA8A12492",
INIT_2D => X"45AAD5400005D7BFFFEFAA800000000000000000000000000000000000000000",
INIT_2E => X"145AAD568B45AAFBFFFEFF7FFD54AAAAAA801EF0000155FFF7FBFDFEFFFD568B",
INIT_2F => X"2155002ABDEBAF7FBFDF55A2AA974AA5D04001EFFFFFD5545557BC21FF080002",
INIT_30 => X"000AA5500174AA0855421FFFFFBEAAAA5D7BEAAAA5D2A82000082E95400A2D54",
INIT_31 => X"BD75FFAAAA80000087BFDF55A2FFE8AAA557FD7410082A800AA557BD74BA0004",
INIT_32 => X"2AAABEF0051400AAA2AAAABFF08003FF55F7FFEABFFF7D57FF455D7FD54105D7",
INIT_33 => X"FD1555FFA2AA800105504001EFFFD140145557BE8BEF000028BEFFFD57FE1000",
INIT_34 => X"0000000000000000000000020005D2E800BA080417400F7FBD75450800174AAF",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000033FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"69844019080000A21A611406840014122A641074155FC28A2024001001801003",
INIT_01 => X"A643D920034004180005E9E3C90360C0041C0181002001602025800008440084",
INIT_02 => X"B7333980808408103F2000F81FC0FEDEAC2161B0B84D0002188011110C018041",
INIT_03 => X"080BA868803F2C020081587008020561E55116B0290000042B71240C800440F8",
INIT_04 => X"42016B0C401F58495C900A4859552A611D9A640F5903B2388004004C08A06008",
INIT_05 => X"16226B107811422A641C08038040007060E0032801E0202000991B708280B501",
INIT_06 => X"B3B8E0FC86142B4142B0000000011114D305824024090A1A143F182000000000",
INIT_07 => X"802102401015610A02C4005000EA019D002482043FCF1C8090C02800C0120886",
INIT_08 => X"20D40A5004003260F9810541494D403D9B98810A0002C601000054B94A006880",
INIT_09 => X"6070000504102805C820C8016C30C250080C0182183804012A0A102200110180",
INIT_0A => X"E000108010230445A800FD865421432121804021C20452880C2D100000022E0C",
INIT_0B => X"C2060014250B9080008306C18360C1B0609C05013065CC042004040808084001",
INIT_0C => X"8582081483ACC15F9C3982081483CCC15F9CBA45505640000A402019003F140F",
INIT_0D => X"F982081483ACC15F9F3982081483CCC15F9FB1962FCB69E08AAAEAEBCDDF7C72",
INIT_0E => X"E3F8E7F5E3AC3620805298B15A3FEBF1CFFF7670ACC3811A28AB57523CDFEBFB",
INIT_0F => X"DC4041D4CF03138DD865103EFEEAC9002BF05800D875E63CC9962FCB52CAA02F",
INIT_10 => X"8DB7BFE25208E8F46A228BF8A757F1B72A8A800B7546DB9F1CA320037F01BD67",
INIT_11 => X"9509EAAE7FD3B749471C48F8A45981CCFAFDBF9464006FD037AEFAE5150016EA",
INIT_12 => X"8802A3AF8E8FB0440CE78773B709641256EC844B8AF92FD7CEDC24A9E181A8A2",
INIT_13 => X"C284601C2864000080113307E4800297D086E00036D2440E0880AAD62BEFF577",
INIT_14 => X"A88DCC2211E44174112840880000060D7030C30B885200D274004008080003C1",
INIT_15 => X"0308003080030800308001840018400400602A01880980037109700C04C44C92",
INIT_16 => X"8340000020301805002D008CD943626111C0D95C20C2030A0030800308003080",
INIT_17 => X"1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B0680834",
INIT_18 => X"B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C",
INIT_19 => X"00000000000041B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1B06C1",
INIT_1A => X"60B22A145DF60B8208209679D701DC2E784601F95163897DF160000000000000",
INIT_1B => X"944A2512AAA8A28A28A2AAAAAA8A28A28A2AAAAAA8A28A28A28A28A28A28A244",
INIT_1C => X"8944A25128944A25128944A25128944A25128944A25128944A25128954AA552A",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8000004A2512",
INIT_1E => X"EAB55FFAA821FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E820BA55000000000000",
INIT_1F => X"16AB55A2D542000A2D5400BA0800021FFFFFFFFFFFFFFBFDFEFAAD142010007B",
INIT_20 => X"80021FFFFFBFDF45A2D56AB45FFFFD54BAFF80001FF002A821FFFFFFFFFEFF7D",
INIT_21 => X"2D140145007BC21FF5D2AAABFFF7D168B45AAD57DFFFFFFFC0010F7842AA10F7",
INIT_22 => X"000002010552E95410AAFBD75FF5D7FEAB5500516AB45A28000010082A975EFA",
INIT_23 => X"5A284155FF5D517FE000004020AA552E80000F7FBC214555003DE10A2FBEAA00",
INIT_24 => X"AA0800154AA0855575FFAAD57FE005D7BD74000804174AA5D00020BA55554214",
INIT_25 => X"0AA490A00000000000000000000000000000000000000000000017400082E954",
INIT_26 => X"AFD7A2D5400001C7BEDB7DEBA4871FFFFFFFFFFFFFFFFDFEFF7FFD74AA552A82",
INIT_27 => X"821FFF7F1F8FC7EBD568B7DB6DF47000AADF400AA080A051FFFFFFFFFEFF7F1F",
INIT_28 => X"1C2000F78A2DA38E38A021C7E3F1F8F55AADB6FB6DFFFBD54AAE38E021FF0824",
INIT_29 => X"8E070281C20925FFBEDB451451C7BC01EF4124ADBC7E3D56AB7DB6DF78FD7EBF",
INIT_2A => X"10E3DE28B6FFE8A101C0E05010412495428AAF1D25EF497FEAB7D145B6FB45AA",
INIT_2B => X"5D0A000BA555F47145BE8A105EF555178E381C0A00092412A87010E3F5C01454",
INIT_2C => X"00000154280024924AA1404174AA0055505EFBEDB7AE385D7FD7438140012482",
INIT_2D => X"EFFFFBD54BA5D2A820AA082A8000000000000000000000000000000000000000",
INIT_2E => X"5FFF7FBFDFEFFFD568B45AAD5400005D7BFFFEFAA80155FFFFFFFFFFFF7FBFDF",
INIT_2F => X"54AAAAAA801EF0000021EFF7D16AB55A2D56ABEFF7FBD5410AAFBC00AA002A95",
INIT_30 => X"68BFFF7FFEAB45AAD140010F7AABFEBAAAAA82145AAD568B45AAFBFFFEFF7FFD",
INIT_31 => X"BE8BFF557BFDF55A2AA974AA5D04001EFFFFFD5545557BC21FF08003FF55AAD1",
INIT_32 => X"2E95400A2D542155002ABDEBAF7FBE8A00552E954100000154AAA2D1421FF007",
INIT_33 => X"D7BD74BA5D0002010552E820AA5D7BD7545F7AA801EF55516AAAA5D2A8200008",
INIT_34 => X"0000000000000000000000174BA0004000AA5500174AA0855421FFFFFBEAAAA5",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000100000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"042200000000000041088001001AA00000000000000000000000500802000003",
INIT_01 => X"200048000024000000000404000000000A22000800000800004A200000000001",
INIT_02 => X"032210008DEF00400060000001C008002489E0F0004037B00010101010000000",
INIT_03 => X"0000010228001000000000000000000024001620280000000000354200004008",
INIT_04 => X"00016200001310090090004840004152C7208802590000388000004C08006000",
INIT_05 => X"1621008008100002641C0803804000702000000000E02000009900000000B100",
INIT_06 => X"0210200C00000000000000000000000080000000000000000003182000000000",
INIT_07 => X"C00D267001B880080700285020020AC98820022802400480405008901100A001",
INIT_08 => X"000000000000106009872048400C4000010D000008000204150A00815A010084",
INIT_09 => X"0000000000000004C80000002C30C200000000021808005800000000000E0E00",
INIT_0A => X"0000000000000000080025860000000080A00020602040800000000000022A04",
INIT_0B => X"C002000000000000000000000000000000000000000000000000000084000760",
INIT_0C => X"385598035D0008A003B05598035D0008A0034078104B41A41000000000031400",
INIT_0D => X"505598035D0008A000B05598035D0008A0004263C0343EDD414004042228DC0D",
INIT_0E => X"0401180DE053A98F6ECC739D8140040231068187C39F5A4F985C008902041124",
INIT_0F => X"227848D4303807FC8CC5508AEAED1BFBD406451B02000E033263C0343CB74050",
INIT_10 => X"00000018A700FCF980CC300318A2420851546B2400000040D8549B5800000010",
INIT_11 => X"40E40511802208D6B30C48F8A8A452210402120A936B0000000004C2A8D64800",
INIT_12 => X"0006362A2B6424287B08286208D6B1427ED430B41402D025082359700181C211",
INIT_13 => X"40000000000000000010030060009C000018440021011821B35254E99AF9E941",
INIT_14 => X"002000044000000000000000000002F0001F00002024B20002000000000002C0",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000040",
INIT_16 => X"00000000000000000000008C8000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"441189B9045D82A69A69803F47E18E0218CC0140400200441920000000000000",
INIT_1B => X"4C261309861861861A69861861861861A69861861861861861861861861861A1",
INIT_1C => X"84C26130984C26130984C26130984C26130984C26130984C261349A4C2613098",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000261309",
INIT_1E => X"820BA55003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A800105D2E8000000000",
INIT_1F => X"FFDFEFF7FFD54BA5D2EA8BFFFF84021FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E",
INIT_20 => X"AE821FFFFFFFFFFFFFFBFDFEFAAD142010007BEAB55FFAABDFFFFFFFFFFFFFFF",
INIT_21 => X"2D542000A2D5400BA08003DFFFFFFFFFFFFF7FBE8B55A2D540010007BEAABAA2",
INIT_22 => X"FFFFFDFEFA2D56AB45AAFBD74AAFFD5420100804021FFFFFFFFFEFF7D16AB55A",
INIT_23 => X"AFF802ABFFFFAE821FFFFFBFDF45A2D56AB45FFFFD54BAFF80001FF002ABDFFF",
INIT_24 => X"45AAD57DFFFFFFFC0010F7842AA10F780155FFF7FBE8B45AAD568BFFF7FBD74B",
INIT_25 => X"000412A8000000000000000000000000000000000000000000002ABFFF7D168B",
INIT_26 => X"DFEFF7FFD74AA552A820AA490A38FFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2A80",
INIT_27 => X"BAFFFFFFFFFFFFF7FBFDFD7EBF1D24AA5D2AADBD7E384071FFFFFFFFFFFFFFFF",
INIT_28 => X"140000007FEFA92A2AA851FFFFFFFFFEFF7F1FAFD7A2D5400001C7BEDB7DEBA4",
INIT_29 => X"F1F8FC7EBD568B7DB6DF47000AADF400AA080A3FFFFFFFBFDFC7E3F5EAB45AAD",
INIT_2A => X"38E021FF0824BDFEFE3F1F8FD7AAD16DB7DBEFBD74AAE3DF400000004021FFF7",
INIT_2B => X"B6DB6FBD7E3F5D04AAFF8A2DBD7E3A0821C7E3F1F8F55AADB6FB6DFFFBD54AAE",
INIT_2C => X"000002DBC7E3D56AB7DB6DF78FD7EBF1C2000F78A2DA38E38A125C7E3F1EAB55",
INIT_2D => X"FFF7FBD54BA552A80010002A8000000000000000000000000000000000000000",
INIT_2E => X"5FFFFFFFFFFFF7FBFDFEFFFFBD54BA5D2A820AA082AA8BFFFFFFFFFFFFFFFFFF",
INIT_2F => X"00005D7BFFFEFAA8028BFFFFFFFDFEFF7FFFFF55A2D5400AA552ABDF55A28015",
INIT_30 => X"FDF55AAD16AB55AAD140010007BFFE10AAAA955FFF7FBFDFEFFFD568B45AAD54",
INIT_31 => X"BC20100800021EFF7D16AB55A2D56ABEFF7FBD5410AAFBC00AA002ABDFEFF7FB",
INIT_32 => X"FBFFFEFF7FFD54AAAAAA801EF00003FFEFA2D56AB45A2D57DFFFFFFFD54AAA2F",
INIT_33 => X"AAA82155AAD568B55FFFFFDF55A2D1400AAF7AABFF45AA8002145AAD568B45AA",
INIT_34 => X"00000000000000000000003FF55AAD168BFFF7FFEAB45AAD140010F7AABFEBAA",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000200000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000003",
INIT_01 => X"A75FF80000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"14088080800008400F655001FFCFF80018FA8044000000000000011000000007",
INIT_03 => X"0000000000000000000000000000000024001660380000000000000000004FF8",
INIT_04 => X"0001E6000053300B00D0005800000000000000407B0004BB830004DC3D01E000",
INIT_05 => X"FEE0000008720043EC3C3D0F87FA19F7E0201C409BE1F10623BB000A100CF300",
INIT_06 => X"06102FFC8E0007C00078008000171175A200096404D9404003FFDBE4744200AA",
INIT_07 => X"482491301000010001DC00000000000000004203FE4005800000008030002000",
INIT_08 => X"20E2008000027FEFF946058180010429000001080AAA010F8000000000000000",
INIT_09 => X"400000120000913FD80000003DF7DE0080010047FBF8000000000800C5408000",
INIT_0A => X"0080000010000400080FFDBE000000400000010000010050600220461003EAFE",
INIT_0B => X"C00600000000801020000000000000010240001721214E000004000000080000",
INIT_0C => X"08020000200000000F30020000200000000F3008001E00000000001803FF14FF",
INIT_0D => X"F0020000200000000F30020000200000000F3040200000020000000026A70C00",
INIT_0E => X"000019B140000800800000020000000030B86000400080000200000000004A58",
INIT_0F => X"AC08000000508001030A0A4001000000000002183E61E6000040200001000000",
INIT_10 => X"0000A56000090100000000001F86C00010080000000000525801000000000014",
INIT_11 => X"0000001716800000803102020000000002BC360020000000000292C010000000",
INIT_12 => X"DF70C08040100000706707600000801000000000000057450000100106060000",
INIT_13 => X"C011001C81080001101F977FE00800000000000040040040002000080506049C",
INIT_14 => X"0000000000000000020020029000000000000000020000000000000000000ADF",
INIT_15 => X"0000000000000000000000000000000000000000000002000200000000000000",
INIT_16 => X"0801810100000000000093ED8000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000401008080",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"930424038000343CF3CF349600704000201120A983400E0104D2040020000000",
INIT_1B => X"190C86432CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB2CB0C30C30C30C30C818",
INIT_1C => X"2190C86432190C86432190C86432190C86432190C86432190C86432190C86432",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8000010C8643",
INIT_1E => X"800105D2EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8201008040000000000",
INIT_1F => X"FFFFFFFFFBD54BA552A8001000003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A",
INIT_20 => X"2E821FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E820BA5500001FFFFFFFFFFFFFF",
INIT_21 => X"7FFD54BA5D2EA8BFFFF843FFFFFFFFFFFFFFFFFFFFEFF7FFD74BA552E801FF00",
INIT_22 => X"FFFFFFFFFFFFBFDFEFFFD542000082EAAB55AAAABDFFFFFFFFFFFFFFFFFDFEFF",
INIT_23 => X"0087BE8B55F784021FFFFFFFFFFFFFFBFDFEFAAD142010007BEAB55FFAA801FF",
INIT_24 => X"FFF7FBE8B55A2D540010007BEAABAA2AE975FFFFFFFFFFFF7FBFDF55AAD14000",
INIT_25 => X"00014000000000000000000000000000000000000000000000003DFFFFFFFFFF",
INIT_26 => X"FFFFFFFBD54AA5D2A80000412ABFFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A82",
INIT_27 => X"021FFFFFFFFFFFFFFFFFFEFF7FBD74BA5D2A800281C0038FFFFFFFFFFFFFFFFF",
INIT_28 => X"FD54BA5D2A801C7142E871FFFFFFFFFFFFFFFFDFEFF7FFD74AA552A820AA490A",
INIT_29 => X"FFFFFFFF7FBFDFD7EBF1D24AA5D2AADBD7E38438FFFFFFFFFFFFFFFBFDFEFFFF",
INIT_2A => X"C7BEDB7DEBA4871FFFFFFFFFEFF7FBF8FD7E3D140010142AAFB7DBEAEBAFFFFF",
INIT_2B => X"E3F1FAF45A2D142010087FEDB55F78A051FFFFFFFFFEFF7F1FAFD7A2D5400001",
INIT_2C => X"000003FFFFFFFBFDFC7E3F5EAB45AAD140000007FEFA92A2AA925FFFFFFFDFEF",
INIT_2D => X"FFFFFFD74AA552A820005D040000000000000000000000000000000000000000",
INIT_2E => X"BFFFFFFFFFFFFFFFFFFFFF7FBD54BA552A80010002ABFFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"54BA5D2A820AA082A821FFFFFFFFFFFFFFBFDFEFF7FFD74AA5D2A800BA550428",
INIT_30 => X"FFFEFF7FBFFFFFF7FBD74BA552A80145552E955FFFFFFFFFFFF7FBFDFEFFFFBD",
INIT_31 => X"ABFFFFFFAEA8BFFFFFFFDFEFF7FFFFF55A2D5400AA552ABDF55A2802ABFFFFFF",
INIT_32 => X"D568B45AAD5400005D7BFFFEFAA80175FFFFFBFDFEFF7FFEAB45AAD1420105D2",
INIT_33 => X"AAA821EFF7FBFDFFFAAD168B55A2D542010007BFDF55F7AE955FFF7FBFDFEFFF",
INIT_34 => X"00000000000000000000003DFEFF7FBFDF55AAD16AB55AAD140010007BFFE10A",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4A302428B824900A128C090A5C1800261500213C005FE812D10420054085A202",
INIT_01 => X"081FFE3440B609703B0427F801A40B8115BC4F655300340288A40D30040E4DD8",
INIT_02 => X"0109095C30C98809800000F9FFFFFFFF149FF1FCA4C0421B182E3490DF145FE4",
INIT_03 => X"1094EC681244819000099486400026523C041660BA000100CC12701015007FF8",
INIT_04 => X"0001E6000053300F01D4587800446194F49020107F0012BBC00202DC3823EA82",
INIT_05 => X"FFF201B228704123FC3C381F87C03DFFF012412A9FE1E01013BF09404050F300",
INIT_06 => X"96F43FFF002004020044041084CB01AD000003761702401000FFDFE050000080",
INIT_07 => X"043C802A821D41412001A0040950AB60014114C3FE4187A009A663A680100B30",
INIT_08 => X"2C01004000047EFFF811A46968004060629A0002208A00000068113205A12034",
INIT_09 => X"0A812D8D5B742D3FF84056383FF7DE0880042107BFF9C45B85101C49A37F4000",
INIT_0A => X"0822189000480406310FFDFE00040009814C089202225412115414601DE3EBFE",
INIT_0B => X"C0281280080180B2948004400220011100841200D001000624000100C002804A",
INIT_0C => X"60694101816002D41A4068C101815004D8158809C86065941840B1014FFF56FF",
INIT_0D => X"0068C101816002D41A40694101815004D815810D42E04A08A80098C024500253",
INIT_0E => X"12682960828F05C96A001B029010134160C8125B0B271802242880A04482418A",
INIT_0F => X"100920C54E8EA256ECF078BA081C10080E05C0B06AA8B12CFD0D42E0441A3000",
INIT_10 => X"4F30A8801406D00290006280320100010362A8A20826A88660D86B202049F115",
INIT_11 => X"2011819E290048A2118EC8140C08064802C0081B0D64040936443306C5514410",
INIT_12 => X"C40A0300600C0A80509F418008804581BA0038005A706680012280506A801060",
INIT_13 => X"C000120080002341881F3FFFF80DCC158092C044600466208CC5091011C322A4",
INIT_14 => X"398C6021569249C4B3007127080806FF917FC30010107688862A28C54518DBFF",
INIT_15 => X"228D9228D9228D9228D99146C9146C84006309044081A001B188300E20806520",
INIT_16 => X"8004000000E07008010003EF80022A51904595123203040D9228D9228D9228D9",
INIT_17 => X"0100401004010040100401004010040100401004010040100401004010044800",
INIT_18 => X"1004010040100401004010040100401004010040100401004010040100401004",
INIT_19 => X"0000000000004010040100401004010040100401004010040100401004010040",
INIT_1A => X"FFBFBFFF7CFE7F9E79E7FFEDDFEFFFBEFFE7DF83F7EFFFFDF7E0000000000000",
INIT_1B => X"FDFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFFD",
INIT_1C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FBFDFEFF7FB",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800003FFFFFF",
INIT_1E => X"8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8001000040000000000",
INIT_1F => X"FFFFFFFFFFD74AA552E80010552EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A",
INIT_20 => X"2ABDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A800105D2EBFFFFFFFFFFFFFFFF",
INIT_21 => X"FFBD54BA552A800100000001FFFFFFFFFFFFFFFFFFFFFFFBD54BA5D2E8201000",
INIT_22 => X"FFFFFFFFFFFFFFFFFFF7FBD74BA5D2E800BA5D00001FFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A552A800BA5D2E821FFFFFFFFFFFFFFFFFFFFF7FBD74AA5D2E820BA5500001FF",
INIT_24 => X"FFFFFFFFFEFF7FFD74BA552E801FF002E975FFFFFFFFFFFFFFFFFFEFF7FBD74A",
INIT_25 => X"00008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA552A8200014003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E80",
INIT_27 => X"BDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2E800005D2ABFFFFFFFFFFFFFFFFFF",
INIT_28 => X"BD54BA552E82028002AB8FFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2A80000412A",
INIT_29 => X"FFFFFFFFFFFFFFEFF7FBD74BA5D2A800281C00001FFFFFFFFFFFFFFFFFFFFF7F",
INIT_2A => X"52A820AA490A071FFFFFFFFFFFFFFFFFFEFF7FBD74AA5D2E800AA5500021FFFF",
INIT_2B => X"FFFFFDFEFF7FFD54BA5D2E80082492E871FFFFFFFFFFFFFFFFDFEFF7FFD74AA5",
INIT_2C => X"0000038FFFFFFFFFFFFFFFBFDFEFFFFFD54BA5D2A801C7142E955FFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8000008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74AA552A820005D043FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"54BA552A80010002ABDFFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2E800005D2EBF",
INIT_30 => X"FFFFFFFFFFDFEFF7FBD74AA552E820BA002AA8BFFFFFFFFFFFFFFFFFFFFF7FBD",
INIT_31 => X"E800BA5D04021FFFFFFFFFFFFFFBFDFEFF7FFD74AA5D2A800BA5504021FFFFFF",
INIT_32 => X"FBFDFEFFFFBD54BA5D2A820AA082A955FFFFFFFFFFFFFFBFDFEFFFFFD54BA552",
INIT_33 => X"52E975FFFFFFFFFEFF7FBFDFFFFFFBD74AA5D2E80000082A955FFFFFFFFFFFF7",
INIT_34 => X"00000000000000000000002ABFFFFFFFFFEFF7FBFFFFFF7FBD74BA552A801455",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"5290F4CDE914905A14A43D33F488243E17122300F55FEB189B343A1140548380",
INIT_01 => X"A94007B259F6A975386262000C344BA9573C6FF57B18A5FB0ABFCD3C2C5F4F0C",
INIT_02 => X"877FE30EB378008D202551040030071869D0040180AC4B685F6E26FAA0810006",
INIT_03 => X"8632CA211E4491D6B5AAD6875AD6AB5A1815600802888808DEA83552954D3000",
INIT_04 => X"24B000808800040439245B221373581F97B0A8D1040F92000F42000047A00E58",
INIT_05 => X"011B2BBA308F023810004700083E220811E9BF2844021B1004045E4249500449",
INIT_06 => X"80A51003AA0200C020088E16A85235722940A817251101010100040D6D0702A2",
INIT_07 => X"5C9ECAB0D247B013B405EAD525FAE48FC2060B880081A26DCD4047EFF9EF0189",
INIT_08 => X"2D0141C0055280100751096B6A40D6F86723E510AA2004803D3275EB2024E814",
INIT_09 => X"04804818CD280100207246A8020000AC0283002004051507A5411C0DA0005048",
INIT_0A => X"2C6898B2950AA65635B00041C23020131A80CFDFF3FE509A907C556828201102",
INIT_0B => X"050F60E220A06880D2A14050A028501428054278142151262CA50343854E506A",
INIT_0C => X"612B3482C0C0078E1F412B1582C090078E1F840A2B0114020104022460002200",
INIT_0D => X"012B1582C0C0078E1F412B3482C090078E1F891C239F8908003099C1ACF06273",
INIT_0E => X"1BA859F213AFC14AA380430060181BA1B0FD16770236A4091621C08055C2C0DB",
INIT_0F => X"B08AA600CA88B143AB11880C280600101F09C030AB28B03C111C239F87082804",
INIT_10 => X"4B61BD8068B92400D0004E30368910E8822A984B0025B0DE6089462660095337",
INIT_11 => X"001AC2173B00E162563454C40804055412D4481128C4CC012A66F30455309600",
INIT_12 => X"50840180A00E1C81900C4190E160589C48082C006A9057CA4385809520F07830",
INIT_13 => X"004416B105036B4180C000800C8C00460848952220592745AC11A544B1BF0068",
INIT_14 => X"512C6A8C4F0008AA800470370000A0004D0000002126F30C902A29C54539C020",
INIT_15 => X"2A81C2A81C2A81C2A81C9540E1540E001400006100003202D040050220103D2A",
INIT_16 => X"22365034A8EA754008004C0214202C50013456520CA09281C2A81C2A81C2A81C",
INIT_17 => X"104411044110441104411044110441104411044110441104411044110445E220",
INIT_18 => X"0401004010040100401004010040100401004411044110441104411044110441",
INIT_19 => X"0003FFFFFFFF9004010040100401004010040100401004010040100401004010",
INIT_1A => X"FFBFAFBEFDFFBBBEFBEFBEFBDFD1FE3EFBD7ADF9B3EFDF7DF7D0512289000000",
INIT_1B => X"FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79EFFC",
INIT_1C => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000FE7F3F",
INIT_1E => X"8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2A8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8201008043FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74AA552E80010552EBFFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E8000055",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD54AA5D2A82000552ABFFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2A800005D2EBDFFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A800105D2EBFFFF",
INIT_24 => X"FFFFFFFFFFFFFFBD54BA5D2E82010002AA8BFFFFFFFFFFFFFFFFFFFFFFFFD54A",
INIT_25 => X"0100004000000000000000000000000000000000000000000000001FFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001008043FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74AA552E800105D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A820001400",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD54AA5D2E800005D2ABFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2A80000412AB8FFFFFFFFFFFFFFFFFFFFFFFFFD54AA5D2A82010552EBDFFFFF",
INIT_2B => X"FFFFFFFFFFFFBD54BA552E80038492EB8FFFFFFFFFFFFFFFFFFFFFFFFBD54AA5",
INIT_2C => X"00000001FFFFFFFFFFFFFFFFFFFFF7FBD54BA552E82028002AA8BFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201000040000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74AA552A820005D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001000043F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD54AA552E8001055003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"A820105D2ABDFFFFFFFFFFFFFFFFFFFFFFFFBD54AA5D2E800005D2EBDFFFFFFF",
INIT_32 => X"FFFFFFFF7FBD54BA552A80010002AA8BFFFFFFFFFFFFFFFFFFFFF7FBD54BA5D2",
INIT_33 => X"02AAABFFFFFFFFFFFFFFFFFFEFF7FBD74BA552E800AA082EA8BFFFFFFFFFFFFF",
INIT_34 => X"0000000000000000000000021FFFFFFFFFFFFFFFFDFEFF7FBD74AA552E820BA0",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"EF20906D902424807BC8241BC81801B97D38AD3C0800103362A6741C80A12A02",
INIT_01 => X"001FFF8409F089003B4422000D80C80106804A7951C5B9D1C828043EA28838F9",
INIT_02 => X"073B8858218C2C50801000F9FFEFF8E72CA7F5FC2E048026496834D84721DFE0",
INIT_03 => X"5886C0201A4001001005080400401420350016E0BB222341C312000014006FF8",
INIT_04 => X"0005EE040057700F40D08078500000D9218020407F0000BB8018A2FC380BEAC2",
INIT_05 => X"FFE0419028700023FCBC385F87C0BFFFE0124002FFE1E0C517FF09111212F300",
INIT_06 => X"16D03FFC96102081020000020489019C430480241202080810FFDFE000000000",
INIT_07 => X"0001160A003475C8100123400E20E1F40F439647FF4807E189A477EF81DF0AF1",
INIT_08 => X"801008000007FEFFFB110140695812CC4188D58A0AAA10803448D0844FB71000",
INIT_09 => X"4201258112D4487FF8001010FFF7DE4000000003BFF8C25818080020017F0F94",
INIT_0A => X"0C024000004A9400000FFDFF50010103134CAFDF03BA18000F39900037C3EBFD",
INIT_0B => X"C02812F00429DC92C40002000100008000105400C00400100000A01800080100",
INIT_0C => X"A1CAF13F214001521001CBF03F21100152100801C17E61841950B1C10FFF57FF",
INIT_0D => X"01CBF03F214001521001CAF13F2110015210088528E00E02C8200A430A424202",
INIT_0E => X"02C86040902AC60BACDF0E02D02001C1C044006D0C94FB94320880603C420B80",
INIT_0F => X"00010AF5052419D196441902801430182800A018D9CA8000648528E00D124802",
INIT_10 => X"4D101808458A5602E000892029110445C19960A00026880C006739000009B003",
INIT_11 => X"1009408021144CB042F880100C0601844068880CE72000013600600332C14000",
INIT_12 => X"F80E02120018390320F050144CB241D0B9023402085020825132C8CB5B404030",
INIT_13 => X"C200400020224000405F7FFFE0008E17C0D240406519400500840A9524EE38A1",
INIT_14 => X"AC810033149249C433200180082A06FF907FC308181204800600000000001BFF",
INIT_15 => X"010C1010C1010C1010C10086080860840063090442A18001B188300C48907120",
INIT_16 => X"0100000000000004002403EFC10302219A41C1443243050C1010C1010C1010C1",
INIT_17 => X"0802008020080200802008020080200802008020080200802008020080200010",
INIT_18 => X"8020080200802008020080200802008020080200802008020080200802008020",
INIT_19 => X"0000000000000080200802008020080200802008020080200802008020080200",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000000000",
INIT_1E => X"8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8001000043FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2A8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA552A8200000043FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A552A8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8201008043FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74AA552E8000055003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2A8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E800000800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA552A8001008043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"52A8200014003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8200008043FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74AA552E820101C003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552E800105D043FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000043F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2A8001008043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"A8200008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA552A8001000043FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74AA552A820005D043FFFFFFFFFFFFFFFFFFFFFFFFFFD74AA552",
INIT_33 => X"5003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA552E8200055043FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003DFFFFFFFFFFFFFFFFFFFFFFFFFD54AA552E800105",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100600007FFF000080108004000800020000840041000080808",
INIT_02 => X"172A00D000EF8210000000F9FFEFF8E7240FF1FC224087B1000639401D005FC0",
INIT_03 => X"0000745C200801000000000400000000340016603A0000004860400014006FFF",
INIT_04 => X"0001E6000053300F00D0007810042140C00000407F0000BB800000DC3801EA00",
INIT_05 => X"FFE0000008700003FC3C380F87C019FFE01240009BE1E00003BF00000000F300",
INIT_06 => X"06103FFC000000000000000004890088010080001202000000FFDFE000000000",
INIT_07 => X"0009B24B043980021000810284204A8001401643FE4007E5501AA00000DC8C30",
INIT_08 => X"0000000000007EFFFB11A56940581280031D61420000B080102040BC5B006120",
INIT_09 => X"020125811254083FF80000003FF7DE0000000003BFF8005800000000017F0000",
INIT_0A => X"0000000000000000000FFDFF4000000AA0354000019C40000128000011C3EBFC",
INIT_0B => X"C000104000000010440000000000000000001000C00000000000000240058000",
INIT_0C => X"4012500021B00880108012500021E00880104809C1666594584031010FFF56FF",
INIT_0D => X"0012500021B00880108012500021E0088010492064206100E81084200048C080",
INIT_0E => X"0410004C840041A0D8005410903804100144800803419043064900C002050184",
INIT_0F => X"020902F60002260D65B361BAA1041018140F02C0000809408D20642053027004",
INIT_10 => X"00020818B06D9802F00030C02060110002C9E8010C00010480B35A0300400041",
INIT_11 => X"20042108603100061516EE800C060228204300166B4060080008240593D00218",
INIT_12 => X"7C02000040206602C10B48110006143B62023C00142800B04400095DFF902030",
INIT_13 => X"C000000000000000001F17FFE000DC1180C7804400044029208301040214AE4C",
INIT_14 => X"008000010012414433000100080806FD107FC300000000000600000000001BFF",
INIT_15 => X"000C1000C1000C1000C100060800608400630104408180012188300C00814080",
INIT_16 => X"0000000000000000000003EF80020201904181003003000C1000C1000C1000C1",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"F30C2416857732AEBAEBFFA55EDCF9822659AE7BE742E6441990000000000000",
INIT_1B => X"3C1E0F07BEFBEFBEF9E79E79E79E79E7BEFBEFBEFBEFBEFBE7BE7BE7BE7BEC98",
INIT_1C => X"83C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F078",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8000001E0F07",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008040000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8001000043FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2A8001000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008040000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100004",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8200008043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8000008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2A8001000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8001000003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008040000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8000008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000043FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8000008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A8000008043FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2A800100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000002015002100000000100000000000000202",
INIT_01 => X"001FFA0000800100200002000000080100004000000020000800041000080808",
INIT_02 => X"1000218000000800000000F9FFEFF8E738FFF1FC20400400000004455A375FE0",
INIT_03 => X"00004000000001000000000400000000340016623A0000004000000014006FFF",
INIT_04 => X"4909E6093253306F82D0007C80000000080E01007F8020BBC00040DC3801EA00",
INIT_05 => X"FFE0000008704503FE3C380F87C019FFF01241009BE1E00203BF80800000F392",
INIT_06 => X"06103FFF9E2086C2086E006604C9019D03108B741202605040FFDFE070400880",
INIT_07 => X"4024057000000100000000000000000001401643FE4007C00000000000CC0830",
INIT_08 => X"0801404000007EFFFF40010000401408000045000000A0801000408000000000",
INIT_09 => X"4A7DF795965C6D3FFC0020003FF7DF01880C618FBFFDD75E00100040437F0000",
INIT_0A => X"0000000000009400000FFDFFC006020000000000019804000028000191C3EBFF",
INIT_0B => X"C02812E0182000F2C48304418220C11160845004D04820000000000000000000",
INIT_0C => X"0002400001000800000002400001000800000801C0786184185031810FFF56FF",
INIT_0D => X"0002400001000800000002400001000800000000202000000800000000080080",
INIT_0E => X"0000000404000000880000001000000001000000000090000008000000040000",
INIT_0F => X"000100C600800001040000040009100000000200200000400000202000020000",
INIT_10 => X"0002000000081001000000000040010000082000000001000001080000000040",
INIT_11 => X"0080000040010000001080001008000000010000210000000008000010400000",
INIT_12 => X"0000030280000000010000010000001020000000000000100400000108000040",
INIT_13 => X"E0120012C1400080291F17FFF0018C11808200400000400000C2000000042000",
INIT_14 => X"00800001001243443B000100880806FD107FC301800000000600000000001BFF",
INIT_15 => X"000C1000C1000C1000C10006080060840077330C4889CC292588300C00804000",
INIT_16 => X"82068C0200000008014023EF80020201904189003003000C1000C1000C1000C1",
INIT_17 => X"110441104411044110441104411044110441104411044110441104451044C820",
INIT_18 => X"1044110441104411044110441104411044110441104411044110441104411044",
INIT_19 => X"FFFFFFFFFFFFC110441104411044110441104411044110441104411044110441",
INIT_1A => X"200A625D144BC2B4D34D7F61432D518B45265EF8278C2015DA080800002FFFFF",
INIT_1B => X"88C4623124924924924924924924924904104104104104104124904124904281",
INIT_1C => X"58AC562B158AC562B158AC562B158AC562B158AC562B158AC56231188C462311",
INIT_1D => X"00000000000000000000000000000000000003FFFFFFFFFFFFFF800002C562B1",
INIT_1E => X"8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8200000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8200000003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"0003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201000043FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"E9264EAB20190CA3BA4997AA9002AE9C001006B0778015CFA17E0811039879C7",
INIT_01 => X"F1FFF9BB1F773C7F9BB07DFFFDD863FC5FFF3FEFFBBF9FFB22FFFBC7B9F30686",
INIT_02 => X"1B33188302E708180F6FFBFFFFCFFFFF9C7FF7FC24350B99082400001D00DFD8",
INIT_03 => X"94A7B2B1450000DCE7366303739CD98C27C57EF57980014F271807E3C9E9CFF8",
INIT_04 => X"6FEBEF5FEC737AFBC6F85FDEB220109E1FEFFFE3FBA7FDFB9BD301DC3FF5F0D2",
INIT_05 => X"FEEDBFDC387F987FEF7C3FAF87FF59F7F5FB7FF59BE1FF980BBBB7FE6D21F3DB",
INIT_06 => X"57902FFDEE9D7DC9D7DF2B263893479DDFAFDFE15213FEFEBFFFFBE1F1D3A333",
INIT_07 => X"10992310605CE10301DE0C1831CB7DF60A244B9BFEE00589DDBCEFEDC1DFA089",
INIT_08 => X"001D8EA111DA7FEFF90F21C8C84D9C0D858FC7020828C18FD18346BBF0000180",
INIT_09 => X"F37DF7B9DF7DCB3FDE89ECC07DF7DF5F985C6BCFFBFA28F99E7EB07F47FFEFAA",
INIT_0A => X"7DCFE1D4077B4D0026FFFFBE7D67D7F3BB79CFFB83BF14EC1E7D5980580BFAFF",
INIT_0B => X"C7D7D51D6F5FDCB935D7AFEBD7F5EBFBF7FEBD66DBFCA3F87501AE7B08060730",
INIT_0C => X"01F45EC0010007E01001F45EC0010007E010084BCD7FF1B61B5C33813FFFFCFF",
INIT_0D => X"01F45EC0010007E01001F45EC0010007E01001BD8020500008001F0100405202",
INIT_0E => X"1EC00040B02007EC09A0E00010001DC0004600400F781429C0080000770001A0",
INIT_0F => X"404B3BFD0402346235408402C08010003C064000E408010081BD802060020000",
INIT_10 => X"0E401A08FE0012040000FC002001360403E434588007200D00F88C84C081C203",
INIT_11 => X"001F01002156040675809145400007B00040091F1190982038406807C868B100",
INIT_12 => X"008320C0403C34000088601604067D00212000007C400082D81009FC08281D00",
INIT_13 => X"F7BFFED3FBFF6A84383F177FF005FFBFF5FA1040076065F730FC08043A903A80",
INIT_14 => X"F589807B7096CD4CF73AC1FC98884FFF19FFC71FEFED7B251E35768E8ED6BFDF",
INIT_15 => X"8C0D78C0D78C0D78C0D7A606BC606B8C56F7730ECCDBDF152199F51EDDCDEBCF",
INIT_16 => X"DFE7DD87FEFF7FF796FFFFFDFFD7E681B867D3683A03A40F78C0D78C0D78C0D7",
INIT_17 => X"BFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEFFBFEFDFD",
INIT_18 => X"FAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFE",
INIT_19 => X"FFFFFFFFFFFFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEBFAFEB",
INIT_1A => X"57AA9ABAD8ACBF0E38E3A89F9E923C2CD990A7D0D2A377F86EDB5C88646FFFFF",
INIT_1B => X"4C261309861861861861861861861861861861861861861861A69A6986186EBC",
INIT_1C => X"84C26130984C26130984C26130984C26130984C26130984C26130984C2613098",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000261309",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100804",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"00080A40000A41248002029000050A088000008242A0004404480002000A1155",
INIT_01 => X"F1FFF1C11F781C129C107DFFFE0860941E81258CA2B71C2220EC1B86E1A00002",
INIT_02 => X"4000002100000014400FF6FFFF0FFFFF8007F1FC211100014200800000887FC0",
INIT_03 => X"1085B0B041000098C63061026318C18404C459757000015F00088BE3C0618FF8",
INIT_04 => X"6FAB975B6470BAF386C87A9CB00000001FEF9F23E3A7BDE79B5101D23FB5C0C2",
INIT_05 => X"F8EDBFD4347F18778E723F2E47FE59C7F5FB7F759B91FB880BA3B6FE2921CBDB",
INIT_06 => X"47000FFC128D5CE8D5CC210638A046889CAB57E8421786B6ACFFE3E181932377",
INIT_07 => X"000000042000000288020C18300320620A80231BFE200181092CE7ED80DFC001",
INIT_08 => X"000C562551D87E8FF90041101042110180004102800008801183468180000141",
INIT_09 => X"137FF7A0FF75813F1C85244071EFBF17D85C738BE3FA08F9DE36B05B07FEEF22",
INIT_0A => X"768EA0C406630D00226FFE3E2D62D6E21259CFDB039E806C02451880400BE0FC",
INIT_0B => X"CC57550D63564D1D2556ADAB56D5AB6AD7EAB962CBD8A3A83101F47E08040510",
INIT_0C => X"01E44A40010007600005E44A4001000760000843C561E5C55C42B9011FFF48FF",
INIT_0D => X"05E44A40010007600005E44A40010007600004BD8020100008001F0100001302",
INIT_0E => X"1EC00000382006EC0820A00010001DC0000208400D781020C008000077000020",
INIT_0F => X"40431BC50402146235400400408010003C064000C400018080BD802020020000",
INIT_10 => X"0E400204FE0010040000FC0000003E0403A424108007200102E888808081C200",
INIT_11 => X"001F0100005E040475808101400007B00000015D111010203840081748482100",
INIT_12 => X"00012040403C34000080201E04047D00202000007C400000F81001FC08080500",
INIT_13 => X"E5ADA4C25ADE72041A3F147FF0018DBBB5FA10400360649310FC08003A903A80",
INIT_14 => X"054880693016DD4C755AC16C1A884FFE18FFD757E7ED7A211E81C09818109E1F",
INIT_15 => X"440C3440C3440C3440C3C2061A2061AD46FF730E5CCBCD55219AB55F0DEFABC7",
INIT_16 => X"5EC71385FC2512E3565BBBF1BAD6F281BC63F1683803C00E3440C3440C3440C3",
INIT_17 => X"B6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6BDE75ED",
INIT_18 => X"6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADA",
INIT_19 => X"FFFFFFFFFFFFAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB6ADAB",
INIT_1A => X"200E5E48710A4200000028150200903950C086D0E28028104A471688747FFFFF",
INIT_1B => X"0080402000000000000000000000000000000000000000020800000000000780",
INIT_1C => X"5028140A05028140A05028140A05028140A05028140A05028140201008040201",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF8000028140A0",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8043FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008043FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"02200AA400180030808802A900002A08001280A08A801044104A1000001818C3",
INIT_01 => X"50A00011460214428114180000882214413D0A71592A01D92213D28005210202",
INIT_02 => X"1444428102100884000AA30200000000C1000401041108404400022220800000",
INIT_03 => X"8C2100804900000C6314A900318C52A40051081000888806108802A141288001",
INIT_04 => X"02000100440408002408008002221000204116A280000F000001400000100010",
INIT_05 => X"0004D44400004D4400000000000000000000005C0000000A0000002C20600000",
INIT_06 => X"4100000120040A0040A00B0090006202940100004000A2020400200888800911",
INIT_07 => X"5002489020420110800244891211440804000810002000081040000000200000",
INIT_08 => X"080542C004CA00000050080202008401842004108AAAA00008912240A1248804",
INIT_09 => X"0000000C0000E400002040500000009202C1002040004400022200020400B062",
INIT_0A => X"58C460540329810002D002000400407020800000004000640800088008280001",
INIT_0B => X"0140000401028008330000800040002002480102010082981500062108020430",
INIT_0C => X"00040A40000000A00000040A40000000A0000040060084104110828030000800",
INIT_0D => X"00040A40000000A00000040A40000000A0000000800010000000000000005000",
INIT_0E => X"00000000A00000040020A000000000000006000000080020C000000000000120",
INIT_0F => X"4040152000000020000004004080000000000000240000000000800020000000",
INIT_10 => X"0000120002000004000000000001220000040410800000090000808080800002",
INIT_11 => X"0000000001420000200001014000000000000900101010200000480008082100",
INIT_12 => X"0001204000000000000820020000200000200000000000028800002000080500",
INIT_13 => X"00933050080C0001900020000000408010000000022000D61028000008000000",
INIT_14 => X"400082D022040000400800081022C0000080000206CB0821082B694D4D294000",
INIT_15 => X"050160501605016050160280B0280B0012000843066021001400040024440245",
INIT_16 => X"0861CD33548542A10209D4100E4040A00002002C004001036050160501605016",
INIT_17 => X"0200802008020080200802008020080200802008020080200802008021081084",
INIT_18 => X"2008020080200802008020080200802008020080200802008020080200802008",
INIT_19 => X"0000000000000020080200802008020080200802008020080200802008020080",
INIT_1A => X"06A0A0F108816B1861863BED822140048D2E5818732C5589A40A0C22E1000000",
INIT_1B => X"80C0603020820820820820820820820820820820820820820820820820820035",
INIT_1C => X"582C160B0582C160B0582C160B0582C160B0582C160B0582C16030180C060301",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800002C160B0",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"000000000000000000000000000000000000000000000003FFFFFFFFC0000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"79964E4BA01DACAB9E659792D00AAE160002829C7FDFEFCEE97C2815039D70C3",
INIT_01 => X"50BFF9AB0775343F9AB01DF80D5821FC0FFF3FEFD1AF9FF1207FFBC7B9720586",
INIT_02 => X"0B33180300E700080F6AAA7BFFC007189C7FF2FC003503980A0000001D00DFD8",
INIT_03 => X"0803B2814D0000C8421A2B03210868AC23403E903900010E271006A148A0C000",
INIT_04 => X"26E1E905CC574828C4F85FC600000016004F77E2F887CDB80BC340DC07D1F000",
INIT_05 => X"FE1DFE4C080F884FE33C078F803F19F011E93ED49BE01F1A03B8972E6D20F049",
INIT_06 => X"57902000DE142D4142D5030010134395D70589415002DA4A17FFF800F0C38111",
INIT_07 => X"00092300601CE00101DE040811D919F402244293FEE00400CCB46BA4C164A088",
INIT_08 => X"08148A4000887FE0000F20C8C80D080D818FC2000000418FD08142BAD0000884",
INIT_09 => X"E204D2154D28AA3FC60888D03C10415A80402847F8002458926A002E457FA0AA",
INIT_0A => X"5587A1540231410006DFFF80540541619968C76980E914E4163D4980100BFA02",
INIT_0B => X"07C7C0140D0B50A8218102C0816040B1225C1506512C83E85500AC3A08040630",
INIT_0C => X"00141EC0000000A01000141EC0000000A01008480D3EB4A24A0C910037FFFC00",
INIT_0D => X"00141EC0000000A01000141EC0000000A0100100800050000000000000405200",
INIT_0E => X"00000040B000010401A0E000000000000046000002080429C0000000000001A0",
INIT_0F => X"40483B590000202000008402C080000000000000240801000100800060000000",
INIT_10 => X"00001A08020002040000000020013600004414588000000D00108484C0800003",
INIT_11 => X"000000002156000220001145400000000040090210909820000068008828B100",
INIT_12 => X"008320C00000000000086016000220000120000000000082D800082000281D00",
INIT_13 => X"32936E43A92F2880B01F37001004B29450580000066021F6303C000408000000",
INIT_14 => X"B481806A62840800C22800B8900042FF0180000ABFEF89250815568A8AD6ABC0",
INIT_15 => X"8D0068D0068D0068D006A68034680300021410028450530014014002D445624D",
INIT_16 => X"89418D13FE7F3FFD8BADB7FC4F4164A00806522C0A40A50268D0068D0068D006",
INIT_17 => X"0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C4B12C9894",
INIT_18 => X"B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C",
INIT_19 => X"FFFFFFFFFFFFC0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0B02C0",
INIT_1A => X"FFBF3F5E7CFC7DFFFFFFD7FADDCFFFBEFFCF1F879DFFFFFDFFEA0C00602FFFFF",
INIT_1B => X"DFEFF7FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBAEBAEBAEBAEBAFFFD",
INIT_1C => X"FDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800003EFF7FB",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"F7AEBEBFFDFFBFBEFBEFFFFFDFF3FC3EFFF7FDFBF76FF7FDFFD0000000000000",
INIT_1B => X"FCFE7F3F9E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79E79EEBD",
INIT_1C => X"9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000FE7F3F",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"129000008004A00804A40000400800020000000C005FEA005800200400050100",
INIT_01 => X"A15FF18019700810180065FFFC0040801E80258CA2951C2200EC0906A0804140",
INIT_02 => X"0000000000000011000550FDFF0FFFFF0007F1FC200000011000000000205FC0",
INIT_03 => X"1084B030000000908428C0024210A30004045060302223490002014280410FF8",
INIT_04 => X"6DA986092050306382C05A1C900000001FAE89016387B2A38B5000D03FA1C0C2",
INIT_05 => X"F8F92B90307F41338E303F0E07FE19C7F1FB7F289B81FB8003A396D20940C3DB",
INIT_06 => X"06000FFC020004C0004C000628800488080003600213001000FFC3E101030222",
INIT_07 => X"000000000000000220000810200220620E00030BFE000181092CE7ED80DF8001",
INIT_08 => X"0000000001107E8FF90001000040100000004102200000801102448100000100",
INIT_09 => X"027DF780DF74013F1C00240071E79F05888C618BA3F800599C101049037E4F40",
INIT_0A => X"240A808004420400202FFC3E002202021259CFDB039E0008024510000023E0FC",
INIT_0B => X"C407500020004C10060204010200810040801060C04821202001A05A00040100",
INIT_0C => X"01E04000010007400001E0400001000740000803C0616184184031010FFF40FF",
INIT_0D => X"01E04000010007400001E04000010007400000BD0020000008001F0100000202",
INIT_0E => X"1EC00000102006E80800000010001DC0000000400D7010000008000077000000",
INIT_0F => X"000308C50402144235400000000010003C064000C000010080BD002000020000",
INIT_10 => X"0E400000FC0010000000FC000000140403A020000007200000E808000001C200",
INIT_11 => X"001F01000014040455808000000007B00000001D010000003840000740400000",
INIT_12 => X"00000000403C34000080001404045D00200000007C400000501001DC08000000",
INIT_13 => X"E004048240426200081F147FF0018C1380DA10400140640100D4080032903A80",
INIT_14 => X"050800A91012494C31004124080886FE187FC301B124F2001600000000001A1F",
INIT_15 => X"000C1000C1000C1000C18006080060840477330C4889CC012188310E08812982",
INIT_16 => X"02061004A820104809402BE1900222019861D1403803800C1000C1000C1000C1",
INIT_17 => X"1004010040100401004010040100401004010040100401004010040100446020",
INIT_18 => X"0040100401004010040100401004010040100401004010040100401004010040",
INIT_19 => X"FFFFFFFFFFFF8100401004010040100401004010040100401004010040100401",
INIT_1A => X"00000000000000000000000000000000000000000000000000001000802FFFFF",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"00000000000000000000000000000000000003007FFFFFFFFFFF800000000000",
INIT_1E => X"8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008000000000000",
INIT_1F => X"FFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E",
INIT_20 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFF",
INIT_21 => X"FFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008",
INIT_22 => X"FFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFF",
INIT_23 => X"A5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFF",
INIT_24 => X"FFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74B",
INIT_25 => X"01008000000000000000000000000000000000000000000000003FFFFFFFFFFF",
INIT_26 => X"FFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E82",
INIT_27 => X"3FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFF",
INIT_28 => X"FD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100800",
INIT_29 => X"FFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_2A => X"D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFF",
INIT_2B => X"FFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5",
INIT_2C => X"000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFF",
INIT_2D => X"FFFFFFD74BA5D2E8201008000000000000000000000000000000000000000000",
INIT_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFF",
INIT_2F => X"74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003F",
INIT_30 => X"FFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD",
INIT_31 => X"E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFF",
INIT_32 => X"FFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2",
INIT_33 => X"8003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E8201008003FFFFFFFFFFFFFFF",
INIT_34 => X"00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFD74BA5D2E820100",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


end;