library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram_plasma is
	port(clk             : in  std_logic;
        address_a       : in  std_logic_vector(31 downto 2);
        enable_a        : in  std_logic;
        wbe_a           : in  std_logic_vector(3 downto 0);
        data_write_a    : in  std_logic_vector(31 downto 0);
        data_read_a     : out std_logic_vector(31 downto 0);

        address_b       : in  std_logic_vector(31 downto 2);
        enable_b        : in  std_logic;
        wbe_b           : in  std_logic_vector(3 downto 0);
        data_write_b    : in  std_logic_vector(31 downto 0);
        data_read_b     : out std_logic_vector(31 downto 0));
end; --entity ram     

architecture ram_plasma of ram_plasma is
signal enable_a_lo       : std_logic;
signal wbe_a_lo          : std_logic_vector(3 downto 0);
signal data_write_a_lo   : std_logic_vector(31 downto 0);
signal data_read_a_lo    : std_logic_vector(31 downto 0);
signal enable_b_lo       : std_logic;
signal wbe_b_lo          : std_logic_vector(3 downto 0);
signal data_read_b_lo    : std_logic_vector(31 downto 0);
signal enable_a_hi       : std_logic;
signal wbe_a_hi          : std_logic_vector(3 downto 0);
signal data_read_a_hi   : std_logic_vector(31 downto 0);
signal enable_b_hi       : std_logic;
signal wbe_b_hi          : std_logic_vector(3 downto 0);
signal data_read_b_hi    : std_logic_vector(31 downto 0);
signal address_a_reg     : std_logic_vector(31 downto 2);
signal address_b_reg     : std_logic_vector(31 downto 2);
signal enable_a_lo_256       : std_logic;
signal wbe_a_lo_256          : std_logic_vector(3 downto 0);
signal data_write_a_lo_256   : std_logic_vector(31 downto 0);
signal data_read_a_lo_256    : std_logic_vector(31 downto 0);
signal enable_b_lo_256       : std_logic;
signal wbe_b_lo_256          : std_logic_vector(3 downto 0);
signal data_read_b_lo_256    : std_logic_vector(31 downto 0);
signal enable_a_hi_256       : std_logic;
signal wbe_a_hi_256          : std_logic_vector(3 downto 0);
signal data_read_a_hi_256   : std_logic_vector(31 downto 0);
signal enable_b_hi_256       : std_logic;
signal wbe_b_hi_256          : std_logic_vector(3 downto 0);
signal data_read_b_hi_256    : std_logic_vector(31 downto 0);
begin
process(clk)
begin
if rising_edge(clk) then
	address_a_reg <= address_a;
	address_b_reg <= address_b;
	end if;
end process;
data_read_a <= data_read_a_lo when (address_a_reg < x"0001000"&"00") else
data_read_a_hi when ((address_a_reg >= x"0001000"&"00") and (address_a_reg < x"0002000"&"00")) else 
data_read_a_lo_256 when ((address_a_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_a_hi_256 when ((address_a_reg >= x"0003000"&"00") and (address_a_reg < x"0004000"&"00"));
data_read_b <= data_read_b_lo when (address_b_reg < x"0001000"&"00") else
data_read_b_hi when ((address_b_reg >= x"0001000"&"00") and (address_b_reg < x"0002000"&"00")) else
data_read_b_lo_256 when ((address_b_reg >= x"0002000"&"00") and (address_a_reg < x"0003000"&"00")) else 
data_read_b_hi_256 when ((address_b_reg >= x"0003000"&"00") and (address_b_reg< x"0004000"&"00"));
enable_a_lo <= enable_a when (address_a < x"0001000"&"00") else '0';
enable_b_lo <= enable_b when (address_b < x"0001000"&"00") else '0';
enable_a_hi <= enable_a when ((address_a >= x"0001000"&"00") and (address_a < x"0002000"&"00")) else '0';
enable_b_hi <= enable_b when ((address_b >= x"0001000"&"00") and (address_b < x"0002000"&"00")) else '0';
enable_a_lo_256 <= enable_a when ((address_a >= x"0002000"&"00") and (address_a < x"0003000"&"00")) else '0';
enable_b_lo_256 <= enable_b when ((address_b >= x"0002000"&"00") and (address_b < x"0003000"&"00")) else '0';
enable_a_hi_256 <= enable_a when ((address_a >= x"0003000"&"00") and (address_a < x"0004000"&"00")) else '0';
enable_b_hi_256 <= enable_b when ((address_b >= x"0003000"&"00") and (address_b < x"0004000"&"00")) else '0';
wbe_a_lo <= wbe_a when  enable_a_lo='1' else x"0";
wbe_a_hi <= wbe_a when  enable_a_hi='1' else x"0";
wbe_b_lo <= wbe_b when  enable_b_lo='1' else x"0";
wbe_b_hi <= wbe_b when  enable_b_hi='1' else x"0";
wbe_a_lo_256 <= wbe_a when  enable_a_lo_256='1' else x"0";
wbe_a_hi_256 <= wbe_a when  enable_a_hi_256='1' else x"0";
wbe_b_lo_256 <= wbe_b when  enable_b_lo_256='1' else x"0";
wbe_b_hi_256 <= wbe_b when  enable_b_hi_256='1' else x"0";



ram_bit_0_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA9918630DD22000000000000128000000400020002106001180000000008003",
INIT_01 => X"80202100005CD2C7B4E6C1E566434955ED29B05AB311C477A91660C2B4D5208F",
INIT_02 => X"11840040D2AC24048604810082640D046B24CC461E01332121AD800087828206",
INIT_03 => X"080029800001E5202400B85242009129400A2A042000F22200808420C4108104",
INIT_04 => X"01FFF3B1EC07842504600200006000844850100838008ED10C280E44011DA811",
INIT_05 => X"3040000004000001A4C949A00000203000010024240D60000C00800242400000",
INIT_06 => X"1E09A28904109024705203C02E348098041390C31050600200958050AA800019",
INIT_07 => X"28AF0779C23B400AF9C0A003557C605D491DA48448900A0208108A05120010E4",
INIT_08 => X"2400008C0010000C00100002008902E8130440D05040C204C2C1312090081370",
INIT_09 => X"0000000000000000000000000000007FE0339694847C449F420A40C368480978",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08451022808200000000000002000000000000010800C000108000000028006",
INIT_01 => X"22402100005000008490005046680400213C00142300E04080F4514BA066C00C",
INIT_02 => X"00000000000020044400010000C28410230CC4480000024000A1800182C12400",
INIT_03 => X"00001000000000000810440001002000802880040000A2020000800004000000",
INIT_04 => X"000DB0B1EC048005006002000028008522200008000004A0000004A002090008",
INIT_05 => X"1480000004000001000800400001210021200090904160000000000909080000",
INIT_06 => X"0008208504104200100000100000901010A1040145448000942100000A808001",
INIT_07 => X"04424205F0124005010C10002000042028092400884080000000020048480048",
INIT_08 => X"A0080004204840040000080A0A200A2A454002080000090A458294C240018200",
INIT_09 => X"0000000000000000000000000000007FE0614546024C1E10064251C088C4057A",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0C0400000682101010101000092D555550554161081447421116AAAAA820012",
INIT_01 => X"0A001DAAA04408028418019800610454A10E00C4000CA262012000C8A0780028",
INIT_02 => X"100400120DC92A5D044335282951264102C1C140091444504A900282D2604003",
INIT_03 => X"82921220A28080400A92560001002012E062020401AE088010808000E4110B00",
INIT_04 => X"100008000200100030000814442D54032820101802A0242A0104843012480048",
INIT_05 => X"14A500A04C448418400080141019210323C258959641002C01550509596D8041",
INIT_06 => X"80A4201F4350564188D54C2852CA5244D2A1011554501081B86100020C10D280",
INIT_07 => X"10405294C0910105021308848045913A20488481D851900022D022084AC9A843",
INIT_08 => X"A14B3D0D0149D2C08680480902A008A21444460200150B9A8D46B4AE500242A9",
INIT_09 => X"0000000000000000000000000000007FF22A53D68064DC5B30EAD404FCF071D0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C100300AE488011001100124C366666619989C84A945469141B33333120002",
INIT_01 => X"0010B50C846428208410028800800004210C0080004802E0558084412581D06C",
INIT_02 => X"1014001A2DC13AA94C09640319D2C44822849441090EA800CA208882C2250108",
INIT_03 => X"3183106A6998924449B054A0100C200804A02200110008904280808005100940",
INIT_04 => X"14000C000000108010002045042B32032829404041B00426108424284A08426A",
INIT_05 => X"0C244E664058850000200011140503090B80449596C8606070CC6109496EC048",
INIT_06 => X"80042815D38052550A05085101C3405452A1010500548530A143160258626300",
INIT_07 => X"024A001480100405020D008060418402A008060020529010218514184A492042",
INIT_08 => X"38D194A5014A7282838524114A19080AC5514649018C09AA954AACA250018A0F",
INIT_09 => X"0000000000000000000000000000007FE350C1460054143016A2C000887031D2",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0CB20AC108100011110000100FC78787806181810800D18195E3C3C3C028006",
INIT_01 => X"081025AA604408128400100081842028A108042040C20260028008C0D4001E2C",
INIT_02 => X"920406000DD1A4110542042879D2002022409101095E64104810200892214103",
INIT_03 => X"87840669E7D0108253B6470800292C1018000000012E28885080601083130802",
INIT_04 => X"40000000000010802080000550370CA52102020207C8240E8380941A3A480026",
INIT_05 => X"0C2151E105000C211022200030214120038000919240406AE3C3212909388059",
INIT_06 => X"00806017E820421400016040008808008481421830255BA49001648258A18424",
INIT_07 => X"8048029480900024440914084041142A20480412804080801784700048488840",
INIT_08 => X"03DB9106014C4282078CE88002083AAE34F30E2B243C299A0D068C8640850008",
INIT_09 => X"0000000000000000000000000000007FED49202102283E622408110054C44518",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"CE88381F030781100000000100D7807F8048181E94A84D60A555C03FC0120006",
INIT_01 => X"083025836054C8D69416D281E46C6D2DA50DA4A0F217E665A82460C84080128C",
INIT_02 => X"918425105D45A411060604228642890040A491071E213031012C8000D7030306",
INIT_03 => X"6860699410016D322448A8D206009113042000042000102A0082501400108001",
INIT_04 => X"55FFF3B1EC0794AD34E02A000040FC8440091018B802AE516C689E45835CB911",
INIT_05 => X"30000C134C5C8880246048952206220929040520221628122C3FA5920220C049",
INIT_06 => X"86ADEA0D46F084351A5B0A506EB686DD148BD0C23D133042100590000000803D",
INIT_07 => X"0AEF157C82B90406B1CD3000653D617FE15C8680B883100328628A1890833CE4",
INIT_08 => X"542D8DA40091A20280520C894A111048030004C0B34352B41A0D190C8001817B",
INIT_09 => X"0000000000000000000000000000017FF07800000EF9FA8F76FC3ED7FDBCFDE9",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4CC0718E26481111111111000D7FF80000FE01E102005601155FFC000000002",
INIT_01 => X"0810258C61440802842102C018619210A10840B00C14B062001008C094001C2C",
INIT_02 => X"120420000090A4110402042000420000088091010002201000200000D0010102",
INIT_03 => X"400010080000000208505481800020D004200004000208000082000000121000",
INIT_04 => X"5400000A10C01088B08168555508028528010000000024204000842102480108",
INIT_05 => X"040008014404088003000604220103210004009594C000024000080959480049",
INIT_06 => X"0084200940205614084100400080800004010000695C48419401100000008000",
INIT_07 => X"800800148090002445090008400100022048049210518081000404004A480840",
INIT_08 => X"A0098004014852138806E8810020080201000E032400299A8D46ACA650850008",
INIT_09 => X"0000000000000000000000000000007FF83BF7F7867CEE7F72EAD507FCFC7CF8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4CC031862648000000000000000000000000000000004000100000000000006",
INIT_01 => X"080025A020440812842112C012099638A10044B009001060000008C014000C2C",
INIT_02 => X"100400020080A4110542042800C2040000809100000220100020000090010002",
INIT_03 => X"4000100800121818484010808040085024200000012C0081D080000000100000",
INIT_04 => X"00000C04120809004010C1000028022009090000000065204001852102CA0428",
INIT_05 => X"C82948000444A41041208215901060020B82100504080000400004A040570400",
INIT_06 => X"0180213F99301D00804044404008800014010800544010411001300250208000",
INIT_07 => X"1008001481941105010910044040100820CA0C81881900018004021002020A51",
INIT_08 => X"00026005010011C102040028081810841500000002000000C060202010010000",
INIT_09 => X"0000000000000000000000000000007FE2000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"D08800000008000000000000000000000000000000800C000100000000000002",
INIT_01 => X"081425A001440802842002C000090410A10800B000140062000001C80080000C",
INIT_02 => X"100400020010A4110542042800420000008011014002200400200000C0010142",
INIT_03 => X"500000080802020000584481840028D204200004000208008080000000301000",
INIT_04 => X"0000004200002040880B00800000020120010000400020005000800102404000",
INIT_05 => X"8400080044040000032006040003250101000191904200805000001909880010",
INIT_06 => X"808400050012420508004840000A804404000001200000409001300000008000",
INIT_07 => X"00080014808000040109100040401000204004009940880110040648C8D92800",
INIT_08 => X"4014190501CA5011880400010200180E010006400200191A0D068C8644210000",
INIT_09 => X"0000000000000000000000000000017FE74B67630200DA6122CCA8C0FCFC7D61",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100204811111111111000000000000000084084C008100000000100002",
INIT_01 => X"000025AAA0440812840112C000609228A10044B00000B060000008C014000C2C",
INIT_02 => X"B20427820090A4110542042801D2046008C00000010264104A302002D2214003",
INIT_03 => X"5000100808000A100850448800202C1014200004012E088050827814C2B20003",
INIT_04 => X"54000C0002081088308028555508020120090000400000A0500010A102014008",
INIT_05 => X"14214803445888001000201120052509090004909250088250000DA909BF8459",
INIT_06 => X"8024488D001242050A404840400A825400004411090100409401300258208000",
INIT_07 => X"020A10948002C4244109100040401108A0016610A942908020040258484B2008",
INIT_08 => X"200000270049E000800404814030080A00200A402200092A158A94CA44210003",
INIT_09 => X"0000000000000000000000000000007FE4234A4E04D5408102225FC4FD58D982",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100264811111111111000000000000000084884C008100000000100002",
INIT_01 => X"081025A360440812840112C000609228A10044B00000B060000808C014000C2C",
INIT_02 => X"100400020010A411054204280152000000801101010220104820000090210102",
INIT_03 => X"4000000800000810004800880020040014200000052C00805080000000100000",
INIT_04 => X"54000C0002081088308028555500028600090000000020004000800102400000",
INIT_05 => X"18214802045C800010202015000642080900050102980800400005B01037C449",
INIT_06 => X"80A0480500200401020008404002025500804001010000411401300A58208000",
INIT_07 => X"024A101080800404020914804040010080400600300310012004041880932800",
INIT_08 => X"400000270081B01000040400423010040100040002001030180C180C00010003",
INIT_09 => X"0000000000000000000000000000007FE771F0778E5016F81494EC15A01C5DA1",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C2880203B0600020202020200000000000400000000004001100000000000006",
INIT_01 => X"0824250C40448882840602C168004100A10180B0B4004064000000C00000000C",
INIT_02 => X"1104001010042411060204000042010000801104540220240024000080010042",
INIT_03 => X"40000888000041002040009302000181042000000000000A8080000000100000",
INIT_04 => X"006AA26948820D258C10C2800000020000010000100000C0402000C103962001",
INIT_05 => X"800008000400000006400C800000000001000000000000004400000000000000",
INIT_06 => X"0401030500000000100000400420000000029800000020401005900000008015",
INIT_07 => X"80840508832D00002489200840184014419604020000000000040000000012B0",
INIT_08 => X"4000040400000010000400080808008014000000120020000000000000850300",
INIT_09 => X"0000000000000000000000000000007FE7394D4E04C1148010440605A158D940",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C88A1F83F000020022002200020000000040004000000480012A000000000002",
INIT_01 => X"081025A00054C8C6940202C06F000801A50080B037810465AA0C60C00000008C",
INIT_02 => X"110400125014A4110746042880428100008411010603302100248000C0030106",
INIT_03 => X"4000018800010400044000DB822095C1142000002000102B8080000000100000",
INIT_04 => X"01F36369D0410025CC5281000040020000011010200000904800008103978000",
INIT_05 => X"E00808004C00000037406E800000000101000000000420004800000000000000",
INIT_06 => X"040D038504000000180002502604008800029C02000000421005B0000000801D",
INIT_07 => X"00000400832EC000820D248065300040019764000000000280048800000012B4",
INIT_08 => X"2400040700000001800400010000000000000000024000000000000000018060",
INIT_09 => X"0000000000000000000000000000007FE701B2B18095005C029A931235189910",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C6CC00100206811133331111580000000000010084084480A320000000100002",
INIT_01 => X"083425A020C40812840552811060DB28A10144A08801F060003809C014000C2C",
INIT_02 => X"114400321014A4110742042803520800408011054102201449240000D4210342",
INIT_03 => X"4800000800016D300048A0880020041014200001832C10A85080020000104400",
INIT_04 => X"559C5DAACECB908DB8EB6AD555400212408901093800EB004C298B010240A800",
INIT_05 => X"0821480244D88004304060910006428909000521229208014C0085B21237C44B",
INIT_06 => X"03ACC805002184000A1002402434028800004002008000411001B0065020801C",
INIT_07 => X"0AA5156880800412B2C9048040306145C04006083083104128040C309092080C",
INIT_08 => X"C00004270091B0008034044140101044020004801A0052341A8D194C82110153",
INIT_09 => X"0000000000000000000000000000017FF83800001EF9FE0F76FC3ED7DDE4E5F8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C088000001600222000000005A0000000040014000000480012A000000000002",
INIT_01 => X"08002500004408028400828000600000A10020A00000A060000000C00000000C",
INIT_02 => X"1084000000002411040204000042000000801100000220000028000081010002",
INIT_03 => X"4000000800000000004000800000000004200000000000000080000000108000",
INIT_04 => X"0001B0E620C72800004202800040020000010000000000004000000102000000",
INIT_05 => X"0000080004000000000000000000000000000000000000004000000000000000",
INIT_06 => X"0000000100000000000000400800000000000000000000401001100000008000",
INIT_07 => X"000000008000000000090000400C000000000400000000000004000000000000",
INIT_08 => X"2000004400000000000400000000000000000000020000000000000000010000",
INIT_09 => X"0000000000000000000000000000007FE07BF7F78E54CEFD36FAFD17FCFC7CF3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08800000060022222222222000000000040000000000400010A000000000002",
INIT_01 => X"08002500004408028400028000000000A10000A000000060000800C00000000C",
INIT_02 => X"1004000000002411040204000042000000A01102160220000020000080010002",
INIT_03 => X"4000298800000000244008800000000004200000000000000080000000100000",
INIT_04 => X"0000001000008564843100000040020000010000000000514000004502000011",
INIT_05 => X"0000080004000000000000000000000000000000000200004000000000000000",
INIT_06 => X"0000000100000020000200400000000000000080000020401001100000008000",
INIT_07 => X"0000000080010000000900004000001000008400000000000804000000000000",
INIT_08 => X"0000000400000000000400000000000000000000020000000000000000010000",
INIT_09 => X"0000000000000000000000000000017FE0000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"05104816EA00C199999999998B82D55555055577C0000675C3816AAAAAB80003",
INIT_01 => X"8014102000081213688B1862C400120ADA22C61962221218A90010E0957F0E0E",
INIT_02 => X"C200BAC50001061C8901300A2C0980A50085C801003641100400A00980206443",
INIT_03 => X"E2D5423CB284889002E20281C02900E8CC00000340A9401040162E6680824001",
INIT_04 => X"FB58CA2929ACA9E021F940410505564001B30303829FBF0A61DAFF19988017A2",
INIT_05 => X"C02C5CB08D408884438B07110220080204209000000028BA6155252000033165",
INIT_06 => X"2420A0A00A840000022800281241080040000208000005E4321254B281295280",
INIT_07 => X"2200000001020208023485003A048820088005000200124342D6311100028200",
INIT_08 => X"91612A8AB000AC00B4C661304000200000110027431500000000001000005485",
INIT_09 => X"0000000000000000000000000000017FE0334A4A0C60F6FB363875D4C538399B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4F74BF57E6E587FFFFFFFFFF92D71999998E665DC000E1D9E8758CCCCCF80000",
INIT_01 => X"2ADE30F033C915094A13393EDEF4B2265284CE4B6F40B85001AE0AB1FA003513",
INIT_02 => X"664123B786736A3991E3A47C1D59727F83855D59A1AC21CA6C30AAA2F8F149E3",
INIT_03 => X"01EF407061DE98DF4182021FC45117E22A0888D2C6F8E0FE6823B275CDE77725",
INIT_04 => X"BB2150ABD272C2B36B5D7FAEEF833D7807BE272701DDBF0600D8FF080FE617A2",
INIT_05 => X"00F1B07EFE79DF5FFF8BFF72DD78043DCFAFDA000117AD7600CF4E60001399BD",
INIT_06 => X"3AFF5F17BF430142FF1415AD12C11700001FF800FCFF5D0421B948FFE3CB1CD7",
INIT_07 => X"77105801B3FDD2780225C3B59F058DB28BFEEC394102168741D8107700029BCB",
INIT_08 => X"A0E66D1FC40024DFE9C023F3F007600088771815600D0020100800010630ECAF",
INIT_09 => X"0000000000000000000000000000017FE00C363180DDE2F82193AAC100343592",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"80900040060040000000000040039E1E1E0F80060E1C067E2F81CF0F0F000003",
INIT_01 => X"82500F0000100211A6110064200002886984501A10005048A99041D0557F0A28",
INIT_02 => X"C0404B0000108804C04211220424A28000C0804940226454001080009001A502",
INIT_03 => X"6078001C3080000000EB02801129001CDC40000100810011D008380302004002",
INIT_04 => X"14CC5F2ABCE128A014BAA8011400FE0280431018808040026081000988000002",
INIT_05 => X"CA0C5C1101DAA0A0038007000206DA400000054342A00210603F31943425E248",
INIT_06 => X"3520A8A040AC0C8020A920A081014C00C208070C000001654B10548004316700",
INIT_07 => X"00005000000104000A360D0295820000000082043609210080661584A1B44430",
INIT_08 => X"90266BAC10A190201046240000001405208005018303969048A41A4C084AD080",
INIT_09 => X"0000000000000000000000000000017FE00917109AA06CA940889D014484C5D9",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"00014020080007FFFFFFFFFF82D7E01FE008005FC000E7E1C1F5F00FF0380003",
INIT_01 => X"0000000000000004108800000000000104220004006A80000000000000000000",
INIT_02 => X"00009440000005400C0000020400000000000000002200000020000940000000",
INIT_03 => X"6040001C3080000000E20280000900000C000000000000000014440010000010",
INIT_04 => X"0031E06403EF80AC801BC19055000E0000030000808000026080000988000002",
INIT_05 => X"00001C1000000000000000000000000000000000000000106003000000060448",
INIT_06 => X"0000000000000000000000100000000000000000000001641063748000048020",
INIT_07 => X"0000000000000000000000002000000000000000000000000046100000000000",
INIT_08 => X"9021104020000000004620000000000000000001030100000000000000000000",
INIT_09 => X"0000000000000000000000000000007FE02EDADE84C87AAA0501480081CC8CB8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"00000000000007FFFFFFFFFF82D7FFE0000FF85FC000E7E1C1F5FFF000380003",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000027C00000180004400007E00000000000000000000",
INIT_03 => X"E7C6867DF780000093E60380000900000C000000000000000000000000000000",
INIT_04 => X"5402305271203D4CC80008550017FE000003000087E2008EE386009BB8190046",
INIT_05 => X"00001DF000000000000000012000008604008000000000F9E3FF000000802803",
INIT_06 => X"0000000000000000000000000000000000000000000003E40000548000000000",
INIT_07 => X"0000000004025200000000000000002008012D000000404007E6700000000000",
INIT_08 => X"33E0040100040C4805EEE00000000000000000230F3F00000000001120000000",
INIT_09 => X"0000000000000000000000000000007FE0402621121D803000120200200848E0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4410801502168D555555555520D7FFFFFF90001F8000057F8D55FFFFFFF00002",
INIT_01 => X"8880BE000439376128C090A2E09240284A30242970600098540084F0017FA04B",
INIT_02 => X"0511481A600817F8800B64437D11428202208800047EF900C80488000085480F",
INIT_03 => X"E7D80EFFF7CC20E513E60BF2044D11000C800040108C0022022B789ECAA60068",
INIT_04 => X"54672E114C020425140002000017FE00050366668780201EE380801FFD140436",
INIT_05 => X"00801FF2120218A12488494149C000200840400200040578E3FF002000170449",
INIT_06 => X"4401A20026C000403008142D00504C00C20E9308545453F43B10568027417811",
INIT_07 => X"1021004806380400821589B43102800083140200010000811FE77000010054A2",
INIT_08 => X"DBF7F9E20001A3C285CFE02200024000A2D500B307BF0020100800000000F056",
INIT_09 => X"0000000000000000000000000000007FE038888C1EF9FE0FF6FC3CD7FDFCFD78",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"6CD0E84501520D555555555524FFFFFFFF90009F8001C17F8055FFFFFFF00000",
INIT_01 => X"0A94BEAFE77D3C314A43D337A45241685290F4CFD22090F85C488C03D57FAC62",
INIT_02 => X"F6157F9A78589FFDD14B756901537001E028C4415900AB14E83DA22A50A5694B",
INIT_03 => X"0827A802001090086000807A1124150890A222023DA002AA52AE78DFEAF6314B",
INIT_04 => X"55F76721460910AD34C028555540006045287676087620400446A00045541AC0",
INIT_05 => X"00A54202485AADB1748AE9510DC4080B28684420220661000000F582022384C9",
INIT_06 => X"54ADCA00000680303A0700FD92A012001036D0C05454D0103B30222A055BFFD5",
INIT_07 => X"1284170066A90561124C8480FA0545630B5480B00288111730018150100258E0",
INIT_08 => X"A817FD23001023D3900105A3409342604044500400800084422111088C6164DF",
INIT_09 => X"0000000000000000000000000000007FE07B77739EF5EEFB76BAFF15E4BCFDF3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"8A99D0720284A800000000006A000000005FFF400C1804002D00000000000002",
INIT_01 => X"A00080000420E3E7BC8241B640909201EF20906F206006E5F4E2B4F0200040CD",
INIT_02 => X"A39050087D451C8190084003FC04B16802C11910167EDC8180382AA20006800C",
INIT_03 => X"E7C02FFFF780000017EE0BA0044D00122CC888D0700CC010020D0094F2A38B73",
INIT_04 => X"019955B0C4038005006002000017FE020003404087818A5FE3980A5FF8000017",
INIT_05 => X"08001FF91300365040888000D01242000282110100900878E3FFF03010124000",
INIT_06 => X"320820000420040000B034B10850100000010004000027F510105680275BFFE8",
INIT_07 => X"000000000000100002134014B008841000000801100108000FF7F40080908000",
INIT_08 => X"1BE000800080100005CFE00000001004A091043B97FF1200000008000002F834",
INIT_09 => X"0000000000000000000000000000007FE0000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010800820001080000840037C00000000000000007E88008380000000040008",
INIT_03 => X"E7C0067FF780000013E603A0000D00000C800000100000000210008001000040",
INIT_04 => X"000CBCB020070000004002000017FE00000340408780000EE380001BF8000006",
INIT_05 => X"00001FF00000000000000000000000000000000000000078E3FFF00000060000",
INIT_06 => X"0000000000000000000000000000000000000000000003F4004C568050200000",
INIT_07 => X"00000000000000000000000004800000000000000000000007E7700000000000",
INIT_08 => X"3BE000400000000005CFE000000000002091002307BF00000000000000000000",
INIT_09 => X"0000000000000000000000000000007FE01D1A18B4B598CC60523ACB39BEBD60",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010000820001080000840037C00028600040000007E88008000000000040008",
INIT_03 => X"E7D8067FF7DC38FD53E623A0000D00000C800000100000000200008000000040",
INIT_04 => X"00000C018C008424042000000017FE00000340408780040EE380041BF8080426",
INIT_05 => X"00001FF000000000000000032224042808040002000004FAE3FFF12020B68010",
INIT_06 => X"00000032FBC009428008000005014C00C2080308000003F40000568000000000",
INIT_07 => X"00A5414910100400B0C0092001022015C00802002102008007E7700001000403",
INIT_08 => X"DBE002201C05A0000DCFE00000002000229108A327BF0230180C100C00000022",
INIT_09 => X"000000000000000000000000000000FFE020272920E9ED0B200C52CF20B83A81",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"85F820440E61E5DDDDDDDDDD81D7FFFFFF8FFE3FDEBCEF7FDFD5FFFFFFF80007",
INIT_01 => X"AA5E3FF033CC1A1BA4993AAC8064328EE9265EAA400ABA7000401AC1DE00573E",
INIT_02 => X"F645FFF78F73EF7DDDE3B57E7C6F72BF89C15D49E0FE675E24302AA9F8D1E5E3",
INIT_03 => X"E7FFD67DF7DE1ADFDBEF578C5479263E7E600053CEFDE25C78BFFE7FDFF77F3F",
INIT_04 => X"FE000C000338529A33843C7FFFBFFF7BAFFF272787FF302EE3D6F03BBE6057EE",
INIT_05 => X"0ED5FDFFF7FBFFFFD889B133FFFFFFFFCFAFDFD7D7FBCFFFE3FF7FFD7DFFFFFF",
INIT_06 => X"38F65C3FFBFF5FD6EFED75ED91C9CF11D688635CE8EB4FE5FBFB7CFDF7FFFFE6",
INIT_07 => X"77525A85B4C017794B3BCFB7DA839D8AAA600FBDFF5BFFC567FE77F7EBFECD03",
INIT_08 => X"B3FFFFFFFDEFFFFFFFEEEFF3F2377C0F29F31F676F3F9DBA9D6EAEBF7E7B7C8F",
INIT_09 => X"000000000000000000000000000000FFE0034B422CD53444E373420BBD2C2CFA",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"11200008002844CCCCCCCCCC80D7FFFFFF8FFE1F5AB4AB7F5ED5FFFFFFEA8015",
INIT_01 => X"080A0E5012800008002029000029049200080A4000142822000002090A800110",
INIT_02 => X"4441D8370DC3416110A004547C8854AB88011100A0FC000A040022202A1000A0",
INIT_03 => X"97EF9671EFDC1ADDDB97570404512A062A000057CA7F0844783D024B19456E38",
INIT_04 => X"FE000C000338529A33843C7FFFBFFDDDAC8E252547F7102E93D6603A3C2056EE",
INIT_05 => X"1611F1FEB2FFF65648209017D9D5B9CECEAA96D6D7798F7D93FF77ED6D7FBFEF",
INIT_06 => X"B0721C3AFBDD5BD7A76D7C05C1CACF55C688231D81804784CF0848A55D7E7BC2",
INIT_07 => X"D35A189424401654452153BC0AC3998AA2200B2BAE5AF54467F873BA6B6FE503",
INIT_08 => X"83FFFF31FD6BEFE677E8EF78FA3E4C8B1D1113474C3F2DAA956AA6BB7AD42E0F",
INIT_09 => X"0000000000000000000000000000007FE03F1110E441278421012A0970222288",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"4128400000606088888888888000000000000000420526004380000000080003",
INIT_01 => X"220A20501184080808802A90006000C202200AA40000A820004A02822A004110",
INIT_02 => X"B24427A5000A440440A21114001A00002288C440A980220A0CA1088828B120A2",
INIT_03 => X"0000000000008000800100041110020C8222220186D182D428827A14E2B25403",
INIT_04 => X"AA000000013042120304142AAA80013881A40303000014000000440000280000",
INIT_05 => X"02B4A005A1A149A7080A1040262094E4E444C2404123C2870000024404803B36",
INIT_06 => X"00523400000B0080050000400000110010352040D4D490005020080D02048002",
INIT_07 => X"41104A01405003310028020040000CA00828019805006CC0500800E220240140",
INIT_08 => X"400000D0E0240C34682002D2B0852621C8444918E80004004000121126310000",
INIT_09 => X"0000000000000000000000000000007FE02064636888C821822C1405C480005B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"A5F0A0540E75C5DDDDDDDDDD81000000000FFE20C60C677EC3D5FFFFFFD80003",
INIT_01 => X"805E1FFFF1C81619E659392E8076B2AE79965E4B402AB858000A0A71FF7FBF3B",
INIT_02 => X"E240FFF78F72EB588DE1A03E016D627D81408809E0FE455E66100001F850C5E1",
INIT_03 => X"E037C67C104E00C793E9038C403806345E4000438F5D604C281FFE7FDFA35F3F",
INIT_04 => X"FE000000013042120304142AAA97FF7A87D72323807E340EE046F41B866813C6",
INIT_05 => X"0A50BC0FF5FBDBBE988131236EBAD6DDC7A78B4141B383FFE0007E541497FF7F",
INIT_06 => X"78D67417992B0592EDA015AC9001010000116000A8AB4BE16BD37C7FF5C57C26",
INIT_07 => X"75100800B0D002380A338E97988008800068051D550176C167FE04F7A0B64941",
INIT_08 => X"9017FFDFE8A4BFFFEDEE03D1B0173405A8A20D37EF00941008040A15263A7481",
INIT_09 => X"0000000000000000000000000000007FE0F480845EF1DE1EFDF8B9DEFDFCFDF8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000222222222225A00000000000140000000800020000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"E000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000007FE03B7F7BFCFDFCEFE37F7E0FFDBCBDF3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_4 : RAMB16_S1_S1
generic map (
INIT_00 => X"60008010001404444444444400D7FFFFFF8FFE1F0810817F0C55FFFFFFE00000",
INIT_01 => X"08800E0FC20105004A40000200128020129000010020000800000030017FA801",
INIT_02 => X"4401D8120D410161100004407D1050EB80011110017C00804A00222200200800",
INIT_03 => X"87EF8671E7DC18DD5386030004410002280888D2492C0080503D004B19452A38",
INIT_04 => X"54000C0002081088308028555517FC40040A242407F7000E83D6201A3C0016E6",
INIT_05 => X"002151FA125AB65040008013D9D4080A0A8A140202100D7883FF75A0203784C9",
INIT_06 => X"60200832FBC40952822D340581C04E00C20C030C000007840B0840A2557A7BC0",
INIT_07 => X"1200100004001440000141B40A83810282000A21220A110427E071100102C403",
INIT_08 => X"03F7FF211C01A3C215C8E5204012400000111007043F00A05028100808402C0F",
INIT_09 => X"0000000000000000000000000000007FE0000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo,               -- Port A enable input
WEA      => wbe_a_lo(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo,               -- Port B enable input
WEB      => wbe_b_lo(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA9918630DD22000000000000128000000400020002106001180000000008003",
INIT_01 => X"80202100005CD2C7B4E6C1E566434955ED29B05AB311C477A91660C2B4D5208F",
INIT_02 => X"11840040D2AC24048604810082640D046B24CC461E01332121AD800087828206",
INIT_03 => X"080029800001E5202400B85242009129400A2A042000F22200808420C4108104",
INIT_04 => X"01FFF3B1EC07842504600200006000844850100838008ED10C280E44011DA811",
INIT_05 => X"3040000004000001A4C949A00000203000010024240D60000C00800242400000",
INIT_06 => X"1E09A28904109024705203C02E348098041390C31050600200958050AA800019",
INIT_07 => X"28AF0779C23B400AF9C0A003557C605D491DA48448900A0208108A05120010E4",
INIT_08 => X"2400008C0010000C00100002008902E8130440D05040C204C2C1312090081370",
INIT_09 => X"0000000000000000000000000000007FE0339694847C449F420A40C368480978",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08451022808200000000000002000000000000010800C000108000000028006",
INIT_01 => X"22402100005000008490005046680400213C00142300E04080F4514BA066C00C",
INIT_02 => X"00000000000020044400010000C28410230CC4480000024000A1800182C12400",
INIT_03 => X"00001000000000000810440001002000802880040000A2020000800004000000",
INIT_04 => X"000DB0B1EC048005006002000028008522200008000004A0000004A002090008",
INIT_05 => X"1480000004000001000800400001210021200090904160000000000909080000",
INIT_06 => X"0008208504104200100000100000901010A1040145448000942100000A808001",
INIT_07 => X"04424205F0124005010C10002000042028092400884080000000020048480048",
INIT_08 => X"A0080004204840040000080A0A200A2A454002080000090A458294C240018200",
INIT_09 => X"0000000000000000000000000000007FE0614546024C1E10064251C088C4057A",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0C0400000682101010101000092D555550554161081447421116AAAAA820012",
INIT_01 => X"0A001DAAA04408028418019800610454A10E00C4000CA262012000C8A0780028",
INIT_02 => X"100400120DC92A5D044335282951264102C1C140091444504A900282D2604003",
INIT_03 => X"82921220A28080400A92560001002012E062020401AE088010808000E4110B00",
INIT_04 => X"100008000200100030000814442D54032820101802A0242A0104843012480048",
INIT_05 => X"14A500A04C448418400080141019210323C258959641002C01550509596D8041",
INIT_06 => X"80A4201F4350564188D54C2852CA5244D2A1011554501081B86100020C10D280",
INIT_07 => X"10405294C0910105021308848045913A20488481D851900022D022084AC9A843",
INIT_08 => X"A14B3D0D0149D2C08680480902A008A21444460200150B9A8D46B4AE500242A9",
INIT_09 => X"0000000000000000000000000000007FF22A53D68064DC5B30EAD404FCF071D0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C100300AE488011001100124C366666619989C84A945469141B33333120002",
INIT_01 => X"0010B50C846428208410028800800004210C0080004802E0558084412581D06C",
INIT_02 => X"1014001A2DC13AA94C09640319D2C44822849441090EA800CA208882C2250108",
INIT_03 => X"3183106A6998924449B054A0100C200804A02200110008904280808005100940",
INIT_04 => X"14000C000000108010002045042B32032829404041B00426108424284A08426A",
INIT_05 => X"0C244E664058850000200011140503090B80449596C8606070CC6109496EC048",
INIT_06 => X"80042815D38052550A05085101C3405452A1010500548530A143160258626300",
INIT_07 => X"024A001480100405020D008060418402A008060020529010218514184A492042",
INIT_08 => X"38D194A5014A7282838524114A19080AC5514649018C09AA954AACA250018A0F",
INIT_09 => X"0000000000000000000000000000007FE350C1460054143016A2C000887031D2",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0CB20AC108100011110000100FC78787806181810800D18195E3C3C3C028006",
INIT_01 => X"081025AA604408128400100081842028A108042040C20260028008C0D4001E2C",
INIT_02 => X"920406000DD1A4110542042879D2002022409101095E64104810200892214103",
INIT_03 => X"87840669E7D0108253B6470800292C1018000000012E28885080601083130802",
INIT_04 => X"40000000000010802080000550370CA52102020207C8240E8380941A3A480026",
INIT_05 => X"0C2151E105000C211022200030214120038000919240406AE3C3212909388059",
INIT_06 => X"00806017E820421400016040008808008481421830255BA49001648258A18424",
INIT_07 => X"8048029480900024440914084041142A20480412804080801784700048488840",
INIT_08 => X"03DB9106014C4282078CE88002083AAE34F30E2B243C299A0D068C8640850008",
INIT_09 => X"0000000000000000000000000000007FED49202102283E622408110054C44518",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"CE88381F030781100000000100D7807F8048181E94A84D60A555C03FC0120006",
INIT_01 => X"083025836054C8D69416D281E46C6D2DA50DA4A0F217E665A82460C84080128C",
INIT_02 => X"918425105D45A411060604228642890040A491071E213031012C8000D7030306",
INIT_03 => X"6860699410016D322448A8D206009113042000042000102A0082501400108001",
INIT_04 => X"55FFF3B1EC0794AD34E02A000040FC8440091018B802AE516C689E45835CB911",
INIT_05 => X"30000C134C5C8880246048952206220929040520221628122C3FA5920220C049",
INIT_06 => X"86ADEA0D46F084351A5B0A506EB686DD148BD0C23D133042100590000000803D",
INIT_07 => X"0AEF157C82B90406B1CD3000653D617FE15C8680B883100328628A1890833CE4",
INIT_08 => X"542D8DA40091A20280520C894A111048030004C0B34352B41A0D190C8001817B",
INIT_09 => X"0000000000000000000000000000017FF07800000EF9FA8F76FC3ED7FDBCFDE9",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4CC0718E26481111111111000D7FF80000FE01E102005601155FFC000000002",
INIT_01 => X"0810258C61440802842102C018619210A10840B00C14B062001008C094001C2C",
INIT_02 => X"120420000090A4110402042000420000088091010002201000200000D0010102",
INIT_03 => X"400010080000000208505481800020D004200004000208000082000000121000",
INIT_04 => X"5400000A10C01088B08168555508028528010000000024204000842102480108",
INIT_05 => X"040008014404088003000604220103210004009594C000024000080959480049",
INIT_06 => X"0084200940205614084100400080800004010000695C48419401100000008000",
INIT_07 => X"800800148090002445090008400100022048049210518081000404004A480840",
INIT_08 => X"A0098004014852138806E8810020080201000E032400299A8D46ACA650850008",
INIT_09 => X"0000000000000000000000000000007FF83BF7F7867CEE7F72EAD507FCFC7CF8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4CC031862648000000000000000000000000000000004000100000000000006",
INIT_01 => X"080025A020440812842112C012099638A10044B009001060000008C014000C2C",
INIT_02 => X"100400020080A4110542042800C2040000809100000220100020000090010002",
INIT_03 => X"4000100800121818484010808040085024200000012C0081D080000000100000",
INIT_04 => X"00000C04120809004010C1000028022009090000000065204001852102CA0428",
INIT_05 => X"C82948000444A41041208215901060020B82100504080000400004A040570400",
INIT_06 => X"0180213F99301D00804044404008800014010800544010411001300250208000",
INIT_07 => X"1008001481941105010910044040100820CA0C81881900018004021002020A51",
INIT_08 => X"00026005010011C102040028081810841500000002000000C060202010010000",
INIT_09 => X"0000000000000000000000000000007FE2000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"D08800000008000000000000000000000000000000800C000100000000000002",
INIT_01 => X"081425A001440802842002C000090410A10800B000140062000001C80080000C",
INIT_02 => X"100400020010A4110542042800420000008011014002200400200000C0010142",
INIT_03 => X"500000080802020000584481840028D204200004000208008080000000301000",
INIT_04 => X"0000004200002040880B00800000020120010000400020005000800102404000",
INIT_05 => X"8400080044040000032006040003250101000191904200805000001909880010",
INIT_06 => X"808400050012420508004840000A804404000001200000409001300000008000",
INIT_07 => X"00080014808000040109100040401000204004009940880110040648C8D92800",
INIT_08 => X"4014190501CA5011880400010200180E010006400200191A0D068C8644210000",
INIT_09 => X"0000000000000000000000000000017FE74B67630200DA6122CCA8C0FCFC7D61",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100204811111111111000000000000000084084C008100000000100002",
INIT_01 => X"000025AAA0440812840112C000609228A10044B00000B060000008C014000C2C",
INIT_02 => X"B20427820090A4110542042801D2046008C00000010264104A302002D2214003",
INIT_03 => X"5000100808000A100850448800202C1014200004012E088050827814C2B20003",
INIT_04 => X"54000C0002081088308028555508020120090000400000A0500010A102014008",
INIT_05 => X"14214803445888001000201120052509090004909250088250000DA909BF8459",
INIT_06 => X"8024488D001242050A404840400A825400004411090100409401300258208000",
INIT_07 => X"020A10948002C4244109100040401108A0016610A942908020040258484B2008",
INIT_08 => X"200000270049E000800404814030080A00200A402200092A158A94CA44210003",
INIT_09 => X"0000000000000000000000000000007FE4234A4E04D5408102225FC4FD58D982",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100264811111111111000000000000000084884C008100000000100002",
INIT_01 => X"081025A360440812840112C000609228A10044B00000B060000808C014000C2C",
INIT_02 => X"100400020010A411054204280152000000801101010220104820000090210102",
INIT_03 => X"4000000800000810004800880020040014200000052C00805080000000100000",
INIT_04 => X"54000C0002081088308028555500028600090000000020004000800102400000",
INIT_05 => X"18214802045C800010202015000642080900050102980800400005B01037C449",
INIT_06 => X"80A0480500200401020008404002025500804001010000411401300A58208000",
INIT_07 => X"024A101080800404020914804040010080400600300310012004041880932800",
INIT_08 => X"400000270081B01000040400423010040100040002001030180C180C00010003",
INIT_09 => X"0000000000000000000000000000007FE771F0778E5016F81494EC15A01C5DA1",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C2880203B0600020202020200000000000400000000004001100000000000006",
INIT_01 => X"0824250C40448882840602C168004100A10180B0B4004064000000C00000000C",
INIT_02 => X"1104001010042411060204000042010000801104540220240024000080010042",
INIT_03 => X"40000888000041002040009302000181042000000000000A8080000000100000",
INIT_04 => X"006AA26948820D258C10C2800000020000010000100000C0402000C103962001",
INIT_05 => X"800008000400000006400C800000000001000000000000004400000000000000",
INIT_06 => X"0401030500000000100000400420000000029800000020401005900000008015",
INIT_07 => X"80840508832D00002489200840184014419604020000000000040000000012B0",
INIT_08 => X"4000040400000010000400080808008014000000120020000000000000850300",
INIT_09 => X"0000000000000000000000000000007FE7394D4E04C1148010440605A158D940",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C88A1F83F000020022002200020000000040004000000480012A000000000002",
INIT_01 => X"081025A00054C8C6940202C06F000801A50080B037810465AA0C60C00000008C",
INIT_02 => X"110400125014A4110746042880428100008411010603302100248000C0030106",
INIT_03 => X"4000018800010400044000DB822095C1142000002000102B8080000000100000",
INIT_04 => X"01F36369D0410025CC5281000040020000011010200000904800008103978000",
INIT_05 => X"E00808004C00000037406E800000000101000000000420004800000000000000",
INIT_06 => X"040D038504000000180002502604008800029C02000000421005B0000000801D",
INIT_07 => X"00000400832EC000820D248065300040019764000000000280048800000012B4",
INIT_08 => X"2400040700000001800400010000000000000000024000000000000000018060",
INIT_09 => X"0000000000000000000000000000007FE701B2B18095005C029A931235189910",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C6CC00100206811133331111580000000000010084084480A320000000100002",
INIT_01 => X"083425A020C40812840552811060DB28A10144A08801F060003809C014000C2C",
INIT_02 => X"114400321014A4110742042803520800408011054102201449240000D4210342",
INIT_03 => X"4800000800016D300048A0880020041014200001832C10A85080020000104400",
INIT_04 => X"559C5DAACECB908DB8EB6AD555400212408901093800EB004C298B010240A800",
INIT_05 => X"0821480244D88004304060910006428909000521229208014C0085B21237C44B",
INIT_06 => X"03ACC805002184000A1002402434028800004002008000411001B0065020801C",
INIT_07 => X"0AA5156880800412B2C9048040306145C04006083083104128040C309092080C",
INIT_08 => X"C00004270091B0008034044140101044020004801A0052341A8D194C82110153",
INIT_09 => X"0000000000000000000000000000017FF83800001EF9FE0F76FC3ED7DDE4E5F8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C088000001600222000000005A0000000040014000000480012A000000000002",
INIT_01 => X"08002500004408028400828000600000A10020A00000A060000000C00000000C",
INIT_02 => X"1084000000002411040204000042000000801100000220000028000081010002",
INIT_03 => X"4000000800000000004000800000000004200000000000000080000000108000",
INIT_04 => X"0001B0E620C72800004202800040020000010000000000004000000102000000",
INIT_05 => X"0000080004000000000000000000000000000000000000004000000000000000",
INIT_06 => X"0000000100000000000000400800000000000000000000401001100000008000",
INIT_07 => X"000000008000000000090000400C000000000400000000000004000000000000",
INIT_08 => X"2000004400000000000400000000000000000000020000000000000000010000",
INIT_09 => X"0000000000000000000000000000007FE07BF7F78E54CEFD36FAFD17FCFC7CF3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08800000060022222222222000000000040000000000400010A000000000002",
INIT_01 => X"08002500004408028400028000000000A10000A000000060000800C00000000C",
INIT_02 => X"1004000000002411040204000042000000A01102160220000020000080010002",
INIT_03 => X"4000298800000000244008800000000004200000000000000080000000100000",
INIT_04 => X"0000001000008564843100000040020000010000000000514000004502000011",
INIT_05 => X"0000080004000000000000000000000000000000000200004000000000000000",
INIT_06 => X"0000000100000020000200400000000000000080000020401001100000008000",
INIT_07 => X"0000000080010000000900004000001000008400000000000804000000000000",
INIT_08 => X"0000000400000000000400000000000000000000020000000000000000010000",
INIT_09 => X"0000000000000000000000000000017FE0000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"05104816EA00C199999999998B82D55555055577C0000675C3816AAAAAB80003",
INIT_01 => X"8014102000081213688B1862C400120ADA22C61962221218A90010E0957F0E0E",
INIT_02 => X"C200BAC50001061C8901300A2C0980A50085C801003641100400A00980206443",
INIT_03 => X"E2D5423CB284889002E20281C02900E8CC00000340A9401040162E6680824001",
INIT_04 => X"FB58CA2929ACA9E021F940410505564001B30303829FBF0A61DAFF19988017A2",
INIT_05 => X"C02C5CB08D408884438B07110220080204209000000028BA6155252000033165",
INIT_06 => X"2420A0A00A840000022800281241080040000208000005E4321254B281295280",
INIT_07 => X"2200000001020208023485003A048820088005000200124342D6311100028200",
INIT_08 => X"91612A8AB000AC00B4C661304000200000110027431500000000001000005485",
INIT_09 => X"0000000000000000000000000000017FE0334A4A0C60F6FB363875D4C538399B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4F74BF57E6E587FFFFFFFFFF92D71999998E665DC000E1D9E8758CCCCCF80000",
INIT_01 => X"2ADE30F033C915094A13393EDEF4B2265284CE4B6F40B85001AE0AB1FA003513",
INIT_02 => X"664123B786736A3991E3A47C1D59727F83855D59A1AC21CA6C30AAA2F8F149E3",
INIT_03 => X"01EF407061DE98DF4182021FC45117E22A0888D2C6F8E0FE6823B275CDE77725",
INIT_04 => X"BB2150ABD272C2B36B5D7FAEEF833D7807BE272701DDBF0600D8FF080FE617A2",
INIT_05 => X"00F1B07EFE79DF5FFF8BFF72DD78043DCFAFDA000117AD7600CF4E60001399BD",
INIT_06 => X"3AFF5F17BF430142FF1415AD12C11700001FF800FCFF5D0421B948FFE3CB1CD7",
INIT_07 => X"77105801B3FDD2780225C3B59F058DB28BFEEC394102168741D8107700029BCB",
INIT_08 => X"A0E66D1FC40024DFE9C023F3F007600088771815600D0020100800010630ECAF",
INIT_09 => X"0000000000000000000000000000017FE00C363180DDE2F82193AAC100343592",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"80900040060040000000000040039E1E1E0F80060E1C067E2F81CF0F0F000003",
INIT_01 => X"82500F0000100211A6110064200002886984501A10005048A99041D0557F0A28",
INIT_02 => X"C0404B0000108804C04211220424A28000C0804940226454001080009001A502",
INIT_03 => X"6078001C3080000000EB02801129001CDC40000100810011D008380302004002",
INIT_04 => X"14CC5F2ABCE128A014BAA8011400FE0280431018808040026081000988000002",
INIT_05 => X"CA0C5C1101DAA0A0038007000206DA400000054342A00210603F31943425E248",
INIT_06 => X"3520A8A040AC0C8020A920A081014C00C208070C000001654B10548004316700",
INIT_07 => X"00005000000104000A360D0295820000000082043609210080661584A1B44430",
INIT_08 => X"90266BAC10A190201046240000001405208005018303969048A41A4C084AD080",
INIT_09 => X"0000000000000000000000000000017FE00917109AA06CA940889D014484C5D9",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"00014020080007FFFFFFFFFF82D7E01FE008005FC000E7E1C1F5F00FF0380003",
INIT_01 => X"0000000000000004108800000000000104220004006A80000000000000000000",
INIT_02 => X"00009440000005400C0000020400000000000000002200000020000940000000",
INIT_03 => X"6040001C3080000000E20280000900000C000000000000000014440010000010",
INIT_04 => X"0031E06403EF80AC801BC19055000E0000030000808000026080000988000002",
INIT_05 => X"00001C1000000000000000000000000000000000000000106003000000060448",
INIT_06 => X"0000000000000000000000100000000000000000000001641063748000048020",
INIT_07 => X"0000000000000000000000002000000000000000000000000046100000000000",
INIT_08 => X"9021104020000000004620000000000000000001030100000000000000000000",
INIT_09 => X"0000000000000000000000000000007FE02EDADE84C87AAA0501480081CC8CB8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"00000000000007FFFFFFFFFF82D7FFE0000FF85FC000E7E1C1F5FFF000380003",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000027C00000180004400007E00000000000000000000",
INIT_03 => X"E7C6867DF780000093E60380000900000C000000000000000000000000000000",
INIT_04 => X"5402305271203D4CC80008550017FE000003000087E2008EE386009BB8190046",
INIT_05 => X"00001DF000000000000000012000008604008000000000F9E3FF000000802803",
INIT_06 => X"0000000000000000000000000000000000000000000003E40000548000000000",
INIT_07 => X"0000000004025200000000000000002008012D000000404007E6700000000000",
INIT_08 => X"33E0040100040C4805EEE00000000000000000230F3F00000000001120000000",
INIT_09 => X"0000000000000000000000000000007FE0402621121D803000120200200848E0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4410801502168D555555555520D7FFFFFF90001F8000057F8D55FFFFFFF00002",
INIT_01 => X"8880BE000439376128C090A2E09240284A30242970600098540084F0017FA04B",
INIT_02 => X"0511481A600817F8800B64437D11428202208800047EF900C80488000085480F",
INIT_03 => X"E7D80EFFF7CC20E513E60BF2044D11000C800040108C0022022B789ECAA60068",
INIT_04 => X"54672E114C020425140002000017FE00050366668780201EE380801FFD140436",
INIT_05 => X"00801FF2120218A12488494149C000200840400200040578E3FF002000170449",
INIT_06 => X"4401A20026C000403008142D00504C00C20E9308545453F43B10568027417811",
INIT_07 => X"1021004806380400821589B43102800083140200010000811FE77000010054A2",
INIT_08 => X"DBF7F9E20001A3C285CFE02200024000A2D500B307BF0020100800000000F056",
INIT_09 => X"0000000000000000000000000000007FE038888C1EF9FE0FF6FC3CD7FDFCFD78",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"6CD0E84501520D555555555524FFFFFFFF90009F8001C17F8055FFFFFFF00000",
INIT_01 => X"0A94BEAFE77D3C314A43D337A45241685290F4CFD22090F85C488C03D57FAC62",
INIT_02 => X"F6157F9A78589FFDD14B756901537001E028C4415900AB14E83DA22A50A5694B",
INIT_03 => X"0827A802001090086000807A1124150890A222023DA002AA52AE78DFEAF6314B",
INIT_04 => X"55F76721460910AD34C028555540006045287676087620400446A00045541AC0",
INIT_05 => X"00A54202485AADB1748AE9510DC4080B28684420220661000000F582022384C9",
INIT_06 => X"54ADCA00000680303A0700FD92A012001036D0C05454D0103B30222A055BFFD5",
INIT_07 => X"1284170066A90561124C8480FA0545630B5480B00288111730018150100258E0",
INIT_08 => X"A817FD23001023D3900105A3409342604044500400800084422111088C6164DF",
INIT_09 => X"0000000000000000000000000000007FE07B77739EF5EEFB76BAFF15E4BCFDF3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"8A99D0720284A800000000006A000000005FFF400C1804002D00000000000002",
INIT_01 => X"A00080000420E3E7BC8241B640909201EF20906F206006E5F4E2B4F0200040CD",
INIT_02 => X"A39050087D451C8190084003FC04B16802C11910167EDC8180382AA20006800C",
INIT_03 => X"E7C02FFFF780000017EE0BA0044D00122CC888D0700CC010020D0094F2A38B73",
INIT_04 => X"019955B0C4038005006002000017FE020003404087818A5FE3980A5FF8000017",
INIT_05 => X"08001FF91300365040888000D01242000282110100900878E3FFF03010124000",
INIT_06 => X"320820000420040000B034B10850100000010004000027F510105680275BFFE8",
INIT_07 => X"000000000000100002134014B008841000000801100108000FF7F40080908000",
INIT_08 => X"1BE000800080100005CFE00000001004A091043B97FF1200000008000002F834",
INIT_09 => X"0000000000000000000000000000007FE0000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010800820001080000840037C00000000000000007E88008380000000040008",
INIT_03 => X"E7C0067FF780000013E603A0000D00000C800000100000000210008001000040",
INIT_04 => X"000CBCB020070000004002000017FE00000340408780000EE380001BF8000006",
INIT_05 => X"00001FF00000000000000000000000000000000000000078E3FFF00000060000",
INIT_06 => X"0000000000000000000000000000000000000000000003F4004C568050200000",
INIT_07 => X"00000000000000000000000004800000000000000000000007E7700000000000",
INIT_08 => X"3BE000400000000005CFE000000000002091002307BF00000000000000000000",
INIT_09 => X"0000000000000000000000000000007FE01D1A18B4B598CC60523ACB39BEBD60",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010000820001080000840037C00028600040000007E88008000000000040008",
INIT_03 => X"E7D8067FF7DC38FD53E623A0000D00000C800000100000000200008000000040",
INIT_04 => X"00000C018C008424042000000017FE00000340408780040EE380041BF8080426",
INIT_05 => X"00001FF000000000000000032224042808040002000004FAE3FFF12020B68010",
INIT_06 => X"00000032FBC009428008000005014C00C2080308000003F40000568000000000",
INIT_07 => X"00A5414910100400B0C0092001022015C00802002102008007E7700001000403",
INIT_08 => X"DBE002201C05A0000DCFE00000002000229108A327BF0230180C100C00000022",
INIT_09 => X"000000000000000000000000000000FFE020272920E9ED0B200C52CF20B83A81",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"85F820440E61E5DDDDDDDDDD81D7FFFFFF8FFE3FDEBCEF7FDFD5FFFFFFF80007",
INIT_01 => X"AA5E3FF033CC1A1BA4993AAC8064328EE9265EAA400ABA7000401AC1DE00573E",
INIT_02 => X"F645FFF78F73EF7DDDE3B57E7C6F72BF89C15D49E0FE675E24302AA9F8D1E5E3",
INIT_03 => X"E7FFD67DF7DE1ADFDBEF578C5479263E7E600053CEFDE25C78BFFE7FDFF77F3F",
INIT_04 => X"FE000C000338529A33843C7FFFBFFF7BAFFF272787FF302EE3D6F03BBE6057EE",
INIT_05 => X"0ED5FDFFF7FBFFFFD889B133FFFFFFFFCFAFDFD7D7FBCFFFE3FF7FFD7DFFFFFF",
INIT_06 => X"38F65C3FFBFF5FD6EFED75ED91C9CF11D688635CE8EB4FE5FBFB7CFDF7FFFFE6",
INIT_07 => X"77525A85B4C017794B3BCFB7DA839D8AAA600FBDFF5BFFC567FE77F7EBFECD03",
INIT_08 => X"B3FFFFFFFDEFFFFFFFEEEFF3F2377C0F29F31F676F3F9DBA9D6EAEBF7E7B7C8F",
INIT_09 => X"000000000000000000000000000000FFE0034B422CD53444E373420BBD2C2CFA",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"11200008002844CCCCCCCCCC80D7FFFFFF8FFE1F5AB4AB7F5ED5FFFFFFEA8015",
INIT_01 => X"080A0E5012800008002029000029049200080A4000142822000002090A800110",
INIT_02 => X"4441D8370DC3416110A004547C8854AB88011100A0FC000A040022202A1000A0",
INIT_03 => X"97EF9671EFDC1ADDDB97570404512A062A000057CA7F0844783D024B19456E38",
INIT_04 => X"FE000C000338529A33843C7FFFBFFDDDAC8E252547F7102E93D6603A3C2056EE",
INIT_05 => X"1611F1FEB2FFF65648209017D9D5B9CECEAA96D6D7798F7D93FF77ED6D7FBFEF",
INIT_06 => X"B0721C3AFBDD5BD7A76D7C05C1CACF55C688231D81804784CF0848A55D7E7BC2",
INIT_07 => X"D35A189424401654452153BC0AC3998AA2200B2BAE5AF54467F873BA6B6FE503",
INIT_08 => X"83FFFF31FD6BEFE677E8EF78FA3E4C8B1D1113474C3F2DAA956AA6BB7AD42E0F",
INIT_09 => X"0000000000000000000000000000007FE03F1110E441278421012A0970222288",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"4128400000606088888888888000000000000000420526004380000000080003",
INIT_01 => X"220A20501184080808802A90006000C202200AA40000A820004A02822A004110",
INIT_02 => X"B24427A5000A440440A21114001A00002288C440A980220A0CA1088828B120A2",
INIT_03 => X"0000000000008000800100041110020C8222220186D182D428827A14E2B25403",
INIT_04 => X"AA000000013042120304142AAA80013881A40303000014000000440000280000",
INIT_05 => X"02B4A005A1A149A7080A1040262094E4E444C2404123C2870000024404803B36",
INIT_06 => X"00523400000B0080050000400000110010352040D4D490005020080D02048002",
INIT_07 => X"41104A01405003310028020040000CA00828019805006CC0500800E220240140",
INIT_08 => X"400000D0E0240C34682002D2B0852621C8444918E80004004000121126310000",
INIT_09 => X"0000000000000000000000000000007FE02064636888C821822C1405C480005B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"A5F0A0540E75C5DDDDDDDDDD81000000000FFE20C60C677EC3D5FFFFFFD80003",
INIT_01 => X"805E1FFFF1C81619E659392E8076B2AE79965E4B402AB858000A0A71FF7FBF3B",
INIT_02 => X"E240FFF78F72EB588DE1A03E016D627D81408809E0FE455E66100001F850C5E1",
INIT_03 => X"E037C67C104E00C793E9038C403806345E4000438F5D604C281FFE7FDFA35F3F",
INIT_04 => X"FE000000013042120304142AAA97FF7A87D72323807E340EE046F41B866813C6",
INIT_05 => X"0A50BC0FF5FBDBBE988131236EBAD6DDC7A78B4141B383FFE0007E541497FF7F",
INIT_06 => X"78D67417992B0592EDA015AC9001010000116000A8AB4BE16BD37C7FF5C57C26",
INIT_07 => X"75100800B0D002380A338E97988008800068051D550176C167FE04F7A0B64941",
INIT_08 => X"9017FFDFE8A4BFFFEDEE03D1B0173405A8A20D37EF00941008040A15263A7481",
INIT_09 => X"0000000000000000000000000000007FE0F480845EF1DE1EFDF8B9DEFDFCFDF8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000222222222225A00000000000140000000800020000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"E000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000007FE03B7F7BFCFDFCEFE37F7E0FFDBCBDF3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_3 : RAMB16_S1_S1
generic map (
INIT_00 => X"60008010001404444444444400D7FFFFFF8FFE1F0810817F0C55FFFFFFE00000",
INIT_01 => X"08800E0FC20105004A40000200128020129000010020000800000030017FA801",
INIT_02 => X"4401D8120D410161100004407D1050EB80011110017C00804A00222200200800",
INIT_03 => X"87EF8671E7DC18DD5386030004410002280888D2492C0080503D004B19452A38",
INIT_04 => X"54000C0002081088308028555517FC40040A242407F7000E83D6201A3C0016E6",
INIT_05 => X"002151FA125AB65040008013D9D4080A0A8A140202100D7883FF75A0203784C9",
INIT_06 => X"60200832FBC40952822D340581C04E00C20C030C000007840B0840A2557A7BC0",
INIT_07 => X"1200100004001440000141B40A83810282000A21220A110427E071100102C403",
INIT_08 => X"03F7FF211C01A3C215C8E5204012400000111007043F00A05028100808402C0F",
INIT_09 => X"0000000000000000000000000000007FE0000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi,               -- Port A enable input
WEA      => wbe_a_hi(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi,               -- Port B enable input
WEB      => wbe_b_hi(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA9918630DD22000000000000128000000400020002106001180000000008003",
INIT_01 => X"80202100005CD2C7B4E6C1E566434955ED29B05AB311C477A91660C2B4D5208F",
INIT_02 => X"11840040D2AC24048604810082640D046B24CC461E01332121AD800087828206",
INIT_03 => X"080029800001E5202400B85242009129400A2A042000F22200808420C4108104",
INIT_04 => X"01FFF3B1EC07842504600200006000844850100838008ED10C280E44011DA811",
INIT_05 => X"3040000004000001A4C949A00000203000010024240D60000C00800242400000",
INIT_06 => X"1E09A28904109024705203C02E348098041390C31050600200958050AA800019",
INIT_07 => X"28AF0779C23B400AF9C0A003557C605D491DA48448900A0208108A05120010E4",
INIT_08 => X"2400008C0010000C00100002008902E8130440D05040C204C2C1312090081370",
INIT_09 => X"0000000000000000000000000000007FE0339694847C449F420A40C368480978",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_lo_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_lo_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08451022808200000000000002000000000000010800C000108000000028006",
INIT_01 => X"22402100005000008490005046680400213C00142300E04080F4514BA066C00C",
INIT_02 => X"00000000000020044400010000C28410230CC4480000024000A1800182C12400",
INIT_03 => X"00001000000000000810440001002000802880040000A2020000800004000000",
INIT_04 => X"000DB0B1EC048005006002000028008522200008000004A0000004A002090008",
INIT_05 => X"1480000004000001000800400001210021200090904160000000000909080000",
INIT_06 => X"0008208504104200100000100000901010A1040145448000942100000A808001",
INIT_07 => X"04424205F0124005010C10002000042028092400884080000000020048480048",
INIT_08 => X"A0080004204840040000080A0A200A2A454002080000090A458294C240018200",
INIT_09 => X"0000000000000000000000000000007FE0614546024C1E10064251C088C4057A",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_lo_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_lo_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0C0400000682101010101000092D555550554161081447421116AAAAA820012",
INIT_01 => X"0A001DAAA04408028418019800610454A10E00C4000CA262012000C8A0780028",
INIT_02 => X"100400120DC92A5D044335282951264102C1C140091444504A900282D2604003",
INIT_03 => X"82921220A28080400A92560001002012E062020401AE088010808000E4110B00",
INIT_04 => X"100008000200100030000814442D54032820101802A0242A0104843012480048",
INIT_05 => X"14A500A04C448418400080141019210323C258959641002C01550509596D8041",
INIT_06 => X"80A4201F4350564188D54C2852CA5244D2A1011554501081B86100020C10D280",
INIT_07 => X"10405294C0910105021308848045913A20488481D851900022D022084AC9A843",
INIT_08 => X"A14B3D0D0149D2C08680480902A008A21444460200150B9A8D46B4AE500242A9",
INIT_09 => X"0000000000000000000000000000007FF22A53D68064DC5B30EAD404FCF071D0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_lo_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_lo_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C100300AE488011001100124C366666619989C84A945469141B33333120002",
INIT_01 => X"0010B50C846428208410028800800004210C0080004802E0558084412581D06C",
INIT_02 => X"1014001A2DC13AA94C09640319D2C44822849441090EA800CA208882C2250108",
INIT_03 => X"3183106A6998924449B054A0100C200804A02200110008904280808005100940",
INIT_04 => X"14000C000000108010002045042B32032829404041B00426108424284A08426A",
INIT_05 => X"0C244E664058850000200011140503090B80449596C8606070CC6109496EC048",
INIT_06 => X"80042815D38052550A05085101C3405452A1010500548530A143160258626300",
INIT_07 => X"024A001480100405020D008060418402A008060020529010218514184A492042",
INIT_08 => X"38D194A5014A7282838524114A19080AC5514649018C09AA954AACA250018A0F",
INIT_09 => X"0000000000000000000000000000007FE350C1460054143016A2C000887031D2",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_lo_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_lo_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0CB20AC108100011110000100FC78787806181810800D18195E3C3C3C028006",
INIT_01 => X"081025AA604408128400100081842028A108042040C20260028008C0D4001E2C",
INIT_02 => X"920406000DD1A4110542042879D2002022409101095E64104810200892214103",
INIT_03 => X"87840669E7D0108253B6470800292C1018000000012E28885080601083130802",
INIT_04 => X"40000000000010802080000550370CA52102020207C8240E8380941A3A480026",
INIT_05 => X"0C2151E105000C211022200030214120038000919240406AE3C3212909388059",
INIT_06 => X"00806017E820421400016040008808008481421830255BA49001648258A18424",
INIT_07 => X"8048029480900024440914084041142A20480412804080801784700048488840",
INIT_08 => X"03DB9106014C4282078CE88002083AAE34F30E2B243C299A0D068C8640850008",
INIT_09 => X"0000000000000000000000000000007FED49202102283E622408110054C44518",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_lo_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_lo_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"CE88381F030781100000000100D7807F8048181E94A84D60A555C03FC0120006",
INIT_01 => X"083025836054C8D69416D281E46C6D2DA50DA4A0F217E665A82460C84080128C",
INIT_02 => X"918425105D45A411060604228642890040A491071E213031012C8000D7030306",
INIT_03 => X"6860699410016D322448A8D206009113042000042000102A0082501400108001",
INIT_04 => X"55FFF3B1EC0794AD34E02A000040FC8440091018B802AE516C689E45835CB911",
INIT_05 => X"30000C134C5C8880246048952206220929040520221628122C3FA5920220C049",
INIT_06 => X"86ADEA0D46F084351A5B0A506EB686DD148BD0C23D133042100590000000803D",
INIT_07 => X"0AEF157C82B90406B1CD3000653D617FE15C8680B883100328628A1890833CE4",
INIT_08 => X"542D8DA40091A20280520C894A111048030004C0B34352B41A0D190C8001817B",
INIT_09 => X"0000000000000000000000000000017FF07800000EF9FA8F76FC3ED7FDBCFDE9",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_lo_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_lo_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4CC0718E26481111111111000D7FF80000FE01E102005601155FFC000000002",
INIT_01 => X"0810258C61440802842102C018619210A10840B00C14B062001008C094001C2C",
INIT_02 => X"120420000090A4110402042000420000088091010002201000200000D0010102",
INIT_03 => X"400010080000000208505481800020D004200004000208000082000000121000",
INIT_04 => X"5400000A10C01088B08168555508028528010000000024204000842102480108",
INIT_05 => X"040008014404088003000604220103210004009594C000024000080959480049",
INIT_06 => X"0084200940205614084100400080800004010000695C48419401100000008000",
INIT_07 => X"800800148090002445090008400100022048049210518081000404004A480840",
INIT_08 => X"A0098004014852138806E8810020080201000E032400299A8D46ACA650850008",
INIT_09 => X"0000000000000000000000000000007FF83BF7F7867CEE7F72EAD507FCFC7CF8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_lo_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_lo_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4CC031862648000000000000000000000000000000004000100000000000006",
INIT_01 => X"080025A020440812842112C012099638A10044B009001060000008C014000C2C",
INIT_02 => X"100400020080A4110542042800C2040000809100000220100020000090010002",
INIT_03 => X"4000100800121818484010808040085024200000012C0081D080000000100000",
INIT_04 => X"00000C04120809004010C1000028022009090000000065204001852102CA0428",
INIT_05 => X"C82948000444A41041208215901060020B82100504080000400004A040570400",
INIT_06 => X"0180213F99301D00804044404008800014010800544010411001300250208000",
INIT_07 => X"1008001481941105010910044040100820CA0C81881900018004021002020A51",
INIT_08 => X"00026005010011C102040028081810841500000002000000C060202010010000",
INIT_09 => X"0000000000000000000000000000007FE2000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_lo_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_lo_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"D08800000008000000000000000000000000000000800C000100000000000002",
INIT_01 => X"081425A001440802842002C000090410A10800B000140062000001C80080000C",
INIT_02 => X"100400020010A4110542042800420000008011014002200400200000C0010142",
INIT_03 => X"500000080802020000584481840028D204200004000208008080000000301000",
INIT_04 => X"0000004200002040880B00800000020120010000400020005000800102404000",
INIT_05 => X"8400080044040000032006040003250101000191904200805000001909880010",
INIT_06 => X"808400050012420508004840000A804404000001200000409001300000008000",
INIT_07 => X"00080014808000040109100040401000204004009940880110040648C8D92800",
INIT_08 => X"4014190501CA5011880400010200180E010006400200191A0D068C8644210000",
INIT_09 => X"0000000000000000000000000000017FE74B67630200DA6122CCA8C0FCFC7D61",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_lo_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_lo_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100204811111111111000000000000000084084C008100000000100002",
INIT_01 => X"000025AAA0440812840112C000609228A10044B00000B060000008C014000C2C",
INIT_02 => X"B20427820090A4110542042801D2046008C00000010264104A302002D2214003",
INIT_03 => X"5000100808000A100850448800202C1014200004012E088050827814C2B20003",
INIT_04 => X"54000C0002081088308028555508020120090000400000A0500010A102014008",
INIT_05 => X"14214803445888001000201120052509090004909250088250000DA909BF8459",
INIT_06 => X"8024488D001242050A404840400A825400004411090100409401300258208000",
INIT_07 => X"020A10948002C4244109100040401108A0016610A942908020040258484B2008",
INIT_08 => X"200000270049E000800404814030080A00200A402200092A158A94CA44210003",
INIT_09 => X"0000000000000000000000000000007FE4234A4E04D5408102225FC4FD58D982",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_lo_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_lo_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100264811111111111000000000000000084884C008100000000100002",
INIT_01 => X"081025A360440812840112C000609228A10044B00000B060000808C014000C2C",
INIT_02 => X"100400020010A411054204280152000000801101010220104820000090210102",
INIT_03 => X"4000000800000810004800880020040014200000052C00805080000000100000",
INIT_04 => X"54000C0002081088308028555500028600090000000020004000800102400000",
INIT_05 => X"18214802045C800010202015000642080900050102980800400005B01037C449",
INIT_06 => X"80A0480500200401020008404002025500804001010000411401300A58208000",
INIT_07 => X"024A101080800404020914804040010080400600300310012004041880932800",
INIT_08 => X"400000270081B01000040400423010040100040002001030180C180C00010003",
INIT_09 => X"0000000000000000000000000000007FE771F0778E5016F81494EC15A01C5DA1",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_lo_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_lo_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C2880203B0600020202020200000000000400000000004001100000000000006",
INIT_01 => X"0824250C40448882840602C168004100A10180B0B4004064000000C00000000C",
INIT_02 => X"1104001010042411060204000042010000801104540220240024000080010042",
INIT_03 => X"40000888000041002040009302000181042000000000000A8080000000100000",
INIT_04 => X"006AA26948820D258C10C2800000020000010000100000C0402000C103962001",
INIT_05 => X"800008000400000006400C800000000001000000000000004400000000000000",
INIT_06 => X"0401030500000000100000400420000000029800000020401005900000008015",
INIT_07 => X"80840508832D00002489200840184014419604020000000000040000000012B0",
INIT_08 => X"4000040400000010000400080808008014000000120020000000000000850300",
INIT_09 => X"0000000000000000000000000000007FE7394D4E04C1148010440605A158D940",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_lo_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_lo_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C88A1F83F000020022002200020000000040004000000480012A000000000002",
INIT_01 => X"081025A00054C8C6940202C06F000801A50080B037810465AA0C60C00000008C",
INIT_02 => X"110400125014A4110746042880428100008411010603302100248000C0030106",
INIT_03 => X"4000018800010400044000DB822095C1142000002000102B8080000000100000",
INIT_04 => X"01F36369D0410025CC5281000040020000011010200000904800008103978000",
INIT_05 => X"E00808004C00000037406E800000000101000000000420004800000000000000",
INIT_06 => X"040D038504000000180002502604008800029C02000000421005B0000000801D",
INIT_07 => X"00000400832EC000820D248065300040019764000000000280048800000012B4",
INIT_08 => X"2400040700000001800400010000000000000000024000000000000000018060",
INIT_09 => X"0000000000000000000000000000007FE701B2B18095005C029A931235189910",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_lo_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_lo_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C6CC00100206811133331111580000000000010084084480A320000000100002",
INIT_01 => X"083425A020C40812840552811060DB28A10144A08801F060003809C014000C2C",
INIT_02 => X"114400321014A4110742042803520800408011054102201449240000D4210342",
INIT_03 => X"4800000800016D300048A0880020041014200001832C10A85080020000104400",
INIT_04 => X"559C5DAACECB908DB8EB6AD555400212408901093800EB004C298B010240A800",
INIT_05 => X"0821480244D88004304060910006428909000521229208014C0085B21237C44B",
INIT_06 => X"03ACC805002184000A1002402434028800004002008000411001B0065020801C",
INIT_07 => X"0AA5156880800412B2C9048040306145C04006083083104128040C309092080C",
INIT_08 => X"C00004270091B0008034044140101044020004801A0052341A8D194C82110153",
INIT_09 => X"0000000000000000000000000000017FF83800001EF9FE0F76FC3ED7DDE4E5F8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_lo_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_lo_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C088000001600222000000005A0000000040014000000480012A000000000002",
INIT_01 => X"08002500004408028400828000600000A10020A00000A060000000C00000000C",
INIT_02 => X"1084000000002411040204000042000000801100000220000028000081010002",
INIT_03 => X"4000000800000000004000800000000004200000000000000080000000108000",
INIT_04 => X"0001B0E620C72800004202800040020000010000000000004000000102000000",
INIT_05 => X"0000080004000000000000000000000000000000000000004000000000000000",
INIT_06 => X"0000000100000000000000400800000000000000000000401001100000008000",
INIT_07 => X"000000008000000000090000400C000000000400000000000004000000000000",
INIT_08 => X"2000004400000000000400000000000000000000020000000000000000010000",
INIT_09 => X"0000000000000000000000000000007FE07BF7F78E54CEFD36FAFD17FCFC7CF3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_lo_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_lo_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08800000060022222222222000000000040000000000400010A000000000002",
INIT_01 => X"08002500004408028400028000000000A10000A000000060000800C00000000C",
INIT_02 => X"1004000000002411040204000042000000A01102160220000020000080010002",
INIT_03 => X"4000298800000000244008800000000004200000000000000080000000100000",
INIT_04 => X"0000001000008564843100000040020000010000000000514000004502000011",
INIT_05 => X"0000080004000000000000000000000000000000000200004000000000000000",
INIT_06 => X"0000000100000020000200400000000000000080000020401001100000008000",
INIT_07 => X"0000000080010000000900004000001000008400000000000804000000000000",
INIT_08 => X"0000000400000000000400000000000000000000020000000000000000010000",
INIT_09 => X"0000000000000000000000000000017FE0000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_lo_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_lo_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"05104816EA00C199999999998B82D55555055577C0000675C3816AAAAAB80003",
INIT_01 => X"8014102000081213688B1862C400120ADA22C61962221218A90010E0957F0E0E",
INIT_02 => X"C200BAC50001061C8901300A2C0980A50085C801003641100400A00980206443",
INIT_03 => X"E2D5423CB284889002E20281C02900E8CC00000340A9401040162E6680824001",
INIT_04 => X"FB58CA2929ACA9E021F940410505564001B30303829FBF0A61DAFF19988017A2",
INIT_05 => X"C02C5CB08D408884438B07110220080204209000000028BA6155252000033165",
INIT_06 => X"2420A0A00A840000022800281241080040000208000005E4321254B281295280",
INIT_07 => X"2200000001020208023485003A048820088005000200124342D6311100028200",
INIT_08 => X"91612A8AB000AC00B4C661304000200000110027431500000000001000005485",
INIT_09 => X"0000000000000000000000000000017FE0334A4A0C60F6FB363875D4C538399B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_lo_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_lo_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4F74BF57E6E587FFFFFFFFFF92D71999998E665DC000E1D9E8758CCCCCF80000",
INIT_01 => X"2ADE30F033C915094A13393EDEF4B2265284CE4B6F40B85001AE0AB1FA003513",
INIT_02 => X"664123B786736A3991E3A47C1D59727F83855D59A1AC21CA6C30AAA2F8F149E3",
INIT_03 => X"01EF407061DE98DF4182021FC45117E22A0888D2C6F8E0FE6823B275CDE77725",
INIT_04 => X"BB2150ABD272C2B36B5D7FAEEF833D7807BE272701DDBF0600D8FF080FE617A2",
INIT_05 => X"00F1B07EFE79DF5FFF8BFF72DD78043DCFAFDA000117AD7600CF4E60001399BD",
INIT_06 => X"3AFF5F17BF430142FF1415AD12C11700001FF800FCFF5D0421B948FFE3CB1CD7",
INIT_07 => X"77105801B3FDD2780225C3B59F058DB28BFEEC394102168741D8107700029BCB",
INIT_08 => X"A0E66D1FC40024DFE9C023F3F007600088771815600D0020100800010630ECAF",
INIT_09 => X"0000000000000000000000000000017FE00C363180DDE2F82193AAC100343592",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_lo_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_lo_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"80900040060040000000000040039E1E1E0F80060E1C067E2F81CF0F0F000003",
INIT_01 => X"82500F0000100211A6110064200002886984501A10005048A99041D0557F0A28",
INIT_02 => X"C0404B0000108804C04211220424A28000C0804940226454001080009001A502",
INIT_03 => X"6078001C3080000000EB02801129001CDC40000100810011D008380302004002",
INIT_04 => X"14CC5F2ABCE128A014BAA8011400FE0280431018808040026081000988000002",
INIT_05 => X"CA0C5C1101DAA0A0038007000206DA400000054342A00210603F31943425E248",
INIT_06 => X"3520A8A040AC0C8020A920A081014C00C208070C000001654B10548004316700",
INIT_07 => X"00005000000104000A360D0295820000000082043609210080661584A1B44430",
INIT_08 => X"90266BAC10A190201046240000001405208005018303969048A41A4C084AD080",
INIT_09 => X"0000000000000000000000000000017FE00917109AA06CA940889D014484C5D9",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_lo_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_lo_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"00014020080007FFFFFFFFFF82D7E01FE008005FC000E7E1C1F5F00FF0380003",
INIT_01 => X"0000000000000004108800000000000104220004006A80000000000000000000",
INIT_02 => X"00009440000005400C0000020400000000000000002200000020000940000000",
INIT_03 => X"6040001C3080000000E20280000900000C000000000000000014440010000010",
INIT_04 => X"0031E06403EF80AC801BC19055000E0000030000808000026080000988000002",
INIT_05 => X"00001C1000000000000000000000000000000000000000106003000000060448",
INIT_06 => X"0000000000000000000000100000000000000000000001641063748000048020",
INIT_07 => X"0000000000000000000000002000000000000000000000000046100000000000",
INIT_08 => X"9021104020000000004620000000000000000001030100000000000000000000",
INIT_09 => X"0000000000000000000000000000007FE02EDADE84C87AAA0501480081CC8CB8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_lo_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_lo_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"00000000000007FFFFFFFFFF82D7FFE0000FF85FC000E7E1C1F5FFF000380003",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000027C00000180004400007E00000000000000000000",
INIT_03 => X"E7C6867DF780000093E60380000900000C000000000000000000000000000000",
INIT_04 => X"5402305271203D4CC80008550017FE000003000087E2008EE386009BB8190046",
INIT_05 => X"00001DF000000000000000012000008604008000000000F9E3FF000000802803",
INIT_06 => X"0000000000000000000000000000000000000000000003E40000548000000000",
INIT_07 => X"0000000004025200000000000000002008012D000000404007E6700000000000",
INIT_08 => X"33E0040100040C4805EEE00000000000000000230F3F00000000001120000000",
INIT_09 => X"0000000000000000000000000000007FE0402621121D803000120200200848E0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_lo_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_lo_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4410801502168D555555555520D7FFFFFF90001F8000057F8D55FFFFFFF00002",
INIT_01 => X"8880BE000439376128C090A2E09240284A30242970600098540084F0017FA04B",
INIT_02 => X"0511481A600817F8800B64437D11428202208800047EF900C80488000085480F",
INIT_03 => X"E7D80EFFF7CC20E513E60BF2044D11000C800040108C0022022B789ECAA60068",
INIT_04 => X"54672E114C020425140002000017FE00050366668780201EE380801FFD140436",
INIT_05 => X"00801FF2120218A12488494149C000200840400200040578E3FF002000170449",
INIT_06 => X"4401A20026C000403008142D00504C00C20E9308545453F43B10568027417811",
INIT_07 => X"1021004806380400821589B43102800083140200010000811FE77000010054A2",
INIT_08 => X"DBF7F9E20001A3C285CFE02200024000A2D500B307BF0020100800000000F056",
INIT_09 => X"0000000000000000000000000000007FE038888C1EF9FE0FF6FC3CD7FDFCFD78",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_lo_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_lo_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"6CD0E84501520D555555555524FFFFFFFF90009F8001C17F8055FFFFFFF00000",
INIT_01 => X"0A94BEAFE77D3C314A43D337A45241685290F4CFD22090F85C488C03D57FAC62",
INIT_02 => X"F6157F9A78589FFDD14B756901537001E028C4415900AB14E83DA22A50A5694B",
INIT_03 => X"0827A802001090086000807A1124150890A222023DA002AA52AE78DFEAF6314B",
INIT_04 => X"55F76721460910AD34C028555540006045287676087620400446A00045541AC0",
INIT_05 => X"00A54202485AADB1748AE9510DC4080B28684420220661000000F582022384C9",
INIT_06 => X"54ADCA00000680303A0700FD92A012001036D0C05454D0103B30222A055BFFD5",
INIT_07 => X"1284170066A90561124C8480FA0545630B5480B00288111730018150100258E0",
INIT_08 => X"A817FD23001023D3900105A3409342604044500400800084422111088C6164DF",
INIT_09 => X"0000000000000000000000000000007FE07B77739EF5EEFB76BAFF15E4BCFDF3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_lo_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_lo_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"8A99D0720284A800000000006A000000005FFF400C1804002D00000000000002",
INIT_01 => X"A00080000420E3E7BC8241B640909201EF20906F206006E5F4E2B4F0200040CD",
INIT_02 => X"A39050087D451C8190084003FC04B16802C11910167EDC8180382AA20006800C",
INIT_03 => X"E7C02FFFF780000017EE0BA0044D00122CC888D0700CC010020D0094F2A38B73",
INIT_04 => X"019955B0C4038005006002000017FE020003404087818A5FE3980A5FF8000017",
INIT_05 => X"08001FF91300365040888000D01242000282110100900878E3FFF03010124000",
INIT_06 => X"320820000420040000B034B10850100000010004000027F510105680275BFFE8",
INIT_07 => X"000000000000100002134014B008841000000801100108000FF7F40080908000",
INIT_08 => X"1BE000800080100005CFE00000001004A091043B97FF1200000008000002F834",
INIT_09 => X"0000000000000000000000000000007FE0000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_lo_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_lo_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010800820001080000840037C00000000000000007E88008380000000040008",
INIT_03 => X"E7C0067FF780000013E603A0000D00000C800000100000000210008001000040",
INIT_04 => X"000CBCB020070000004002000017FE00000340408780000EE380001BF8000006",
INIT_05 => X"00001FF00000000000000000000000000000000000000078E3FFF00000060000",
INIT_06 => X"0000000000000000000000000000000000000000000003F4004C568050200000",
INIT_07 => X"00000000000000000000000004800000000000000000000007E7700000000000",
INIT_08 => X"3BE000400000000005CFE000000000002091002307BF00000000000000000000",
INIT_09 => X"0000000000000000000000000000007FE01D1A18B4B598CC60523ACB39BEBD60",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_lo_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_lo_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010000820001080000840037C00028600040000007E88008000000000040008",
INIT_03 => X"E7D8067FF7DC38FD53E623A0000D00000C800000100000000200008000000040",
INIT_04 => X"00000C018C008424042000000017FE00000340408780040EE380041BF8080426",
INIT_05 => X"00001FF000000000000000032224042808040002000004FAE3FFF12020B68010",
INIT_06 => X"00000032FBC009428008000005014C00C2080308000003F40000568000000000",
INIT_07 => X"00A5414910100400B0C0092001022015C00802002102008007E7700001000403",
INIT_08 => X"DBE002201C05A0000DCFE00000002000229108A327BF0230180C100C00000022",
INIT_09 => X"000000000000000000000000000000FFE020272920E9ED0B200C52CF20B83A81",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_lo_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_lo_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"85F820440E61E5DDDDDDDDDD81D7FFFFFF8FFE3FDEBCEF7FDFD5FFFFFFF80007",
INIT_01 => X"AA5E3FF033CC1A1BA4993AAC8064328EE9265EAA400ABA7000401AC1DE00573E",
INIT_02 => X"F645FFF78F73EF7DDDE3B57E7C6F72BF89C15D49E0FE675E24302AA9F8D1E5E3",
INIT_03 => X"E7FFD67DF7DE1ADFDBEF578C5479263E7E600053CEFDE25C78BFFE7FDFF77F3F",
INIT_04 => X"FE000C000338529A33843C7FFFBFFF7BAFFF272787FF302EE3D6F03BBE6057EE",
INIT_05 => X"0ED5FDFFF7FBFFFFD889B133FFFFFFFFCFAFDFD7D7FBCFFFE3FF7FFD7DFFFFFF",
INIT_06 => X"38F65C3FFBFF5FD6EFED75ED91C9CF11D688635CE8EB4FE5FBFB7CFDF7FFFFE6",
INIT_07 => X"77525A85B4C017794B3BCFB7DA839D8AAA600FBDFF5BFFC567FE77F7EBFECD03",
INIT_08 => X"B3FFFFFFFDEFFFFFFFEEEFF3F2377C0F29F31F676F3F9DBA9D6EAEBF7E7B7C8F",
INIT_09 => X"000000000000000000000000000000FFE0034B422CD53444E373420BBD2C2CFA",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_lo_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_lo_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"11200008002844CCCCCCCCCC80D7FFFFFF8FFE1F5AB4AB7F5ED5FFFFFFEA8015",
INIT_01 => X"080A0E5012800008002029000029049200080A4000142822000002090A800110",
INIT_02 => X"4441D8370DC3416110A004547C8854AB88011100A0FC000A040022202A1000A0",
INIT_03 => X"97EF9671EFDC1ADDDB97570404512A062A000057CA7F0844783D024B19456E38",
INIT_04 => X"FE000C000338529A33843C7FFFBFFDDDAC8E252547F7102E93D6603A3C2056EE",
INIT_05 => X"1611F1FEB2FFF65648209017D9D5B9CECEAA96D6D7798F7D93FF77ED6D7FBFEF",
INIT_06 => X"B0721C3AFBDD5BD7A76D7C05C1CACF55C688231D81804784CF0848A55D7E7BC2",
INIT_07 => X"D35A189424401654452153BC0AC3998AA2200B2BAE5AF54467F873BA6B6FE503",
INIT_08 => X"83FFFF31FD6BEFE677E8EF78FA3E4C8B1D1113474C3F2DAA956AA6BB7AD42E0F",
INIT_09 => X"0000000000000000000000000000007FE03F1110E441278421012A0970222288",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_lo_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_lo_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"4128400000606088888888888000000000000000420526004380000000080003",
INIT_01 => X"220A20501184080808802A90006000C202200AA40000A820004A02822A004110",
INIT_02 => X"B24427A5000A440440A21114001A00002288C440A980220A0CA1088828B120A2",
INIT_03 => X"0000000000008000800100041110020C8222220186D182D428827A14E2B25403",
INIT_04 => X"AA000000013042120304142AAA80013881A40303000014000000440000280000",
INIT_05 => X"02B4A005A1A149A7080A1040262094E4E444C2404123C2870000024404803B36",
INIT_06 => X"00523400000B0080050000400000110010352040D4D490005020080D02048002",
INIT_07 => X"41104A01405003310028020040000CA00828019805006CC0500800E220240140",
INIT_08 => X"400000D0E0240C34682002D2B0852621C8444918E80004004000121126310000",
INIT_09 => X"0000000000000000000000000000007FE02064636888C821822C1405C480005B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_lo_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_lo_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"A5F0A0540E75C5DDDDDDDDDD81000000000FFE20C60C677EC3D5FFFFFFD80003",
INIT_01 => X"805E1FFFF1C81619E659392E8076B2AE79965E4B402AB858000A0A71FF7FBF3B",
INIT_02 => X"E240FFF78F72EB588DE1A03E016D627D81408809E0FE455E66100001F850C5E1",
INIT_03 => X"E037C67C104E00C793E9038C403806345E4000438F5D604C281FFE7FDFA35F3F",
INIT_04 => X"FE000000013042120304142AAA97FF7A87D72323807E340EE046F41B866813C6",
INIT_05 => X"0A50BC0FF5FBDBBE988131236EBAD6DDC7A78B4141B383FFE0007E541497FF7F",
INIT_06 => X"78D67417992B0592EDA015AC9001010000116000A8AB4BE16BD37C7FF5C57C26",
INIT_07 => X"75100800B0D002380A338E97988008800068051D550176C167FE04F7A0B64941",
INIT_08 => X"9017FFDFE8A4BFFFEDEE03D1B0173405A8A20D37EF00941008040A15263A7481",
INIT_09 => X"0000000000000000000000000000007FE0F480845EF1DE1EFDF8B9DEFDFCFDF8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_lo_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_lo_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000222222222225A00000000000140000000800020000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"E000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000007FE03B7F7BFCFDFCEFE37F7E0FFDBCBDF3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_lo_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_lo_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_2 : RAMB16_S1_S1
generic map (
INIT_00 => X"60008010001404444444444400D7FFFFFF8FFE1F0810817F0C55FFFFFFE00000",
INIT_01 => X"08800E0FC20105004A40000200128020129000010020000800000030017FA801",
INIT_02 => X"4401D8120D410161100004407D1050EB80011110017C00804A00222200200800",
INIT_03 => X"87EF8671E7DC18DD5386030004410002280888D2492C0080503D004B19452A38",
INIT_04 => X"54000C0002081088308028555517FC40040A242407F7000E83D6201A3C0016E6",
INIT_05 => X"002151FA125AB65040008013D9D4080A0A8A140202100D7883FF75A0203784C9",
INIT_06 => X"60200832FBC40952822D340581C04E00C20C030C000007840B0840A2557A7BC0",
INIT_07 => X"1200100004001440000141B40A83810282000A21220A110427E071100102C403",
INIT_08 => X"03F7FF211C01A3C215C8E5204012400000111007043F00A05028100808402C0F",
INIT_09 => X"0000000000000000000000000000007FE0000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_lo_256,               -- Port A enable input
WEA      => wbe_a_lo_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_lo_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_lo_256,               -- Port B enable input
WEB      => wbe_b_lo_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_lo_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_0_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"DA9918630DD22000000000000128000000400020002106001180000000008003",
INIT_01 => X"80202100005CD2C7B4E6C1E566434955ED29B05AB311C477A91660C2B4D5208F",
INIT_02 => X"11840040D2AC24048604810082640D046B24CC461E01332121AD800087828206",
INIT_03 => X"080029800001E5202400B85242009129400A2A042000F22200808420C4108104",
INIT_04 => X"01FFF3B1EC07842504600200006000844850100838008ED10C280E44011DA811",
INIT_05 => X"3040000004000001A4C949A00000203000010024240D60000C00800242400000",
INIT_06 => X"1E09A28904109024705203C02E348098041390C31050600200958050AA800019",
INIT_07 => X"28AF0779C23B400AF9C0A003557C605D491DA48448900A0208108A05120010E4",
INIT_08 => X"2400008C0010000C00100002008902E8130440D05040C204C2C1312090081370",
INIT_09 => X"0000000000000000000000000000007FE0339694847C449F420A40C368480978",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(0),        -- Port A data input
DOA(0)   => data_read_a_hi_256(0),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(0),        -- Port B data input
DOB(0)   => data_read_b_hi_256(0),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_1_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08451022808200000000000002000000000000010800C000108000000028006",
INIT_01 => X"22402100005000008490005046680400213C00142300E04080F4514BA066C00C",
INIT_02 => X"00000000000020044400010000C28410230CC4480000024000A1800182C12400",
INIT_03 => X"00001000000000000810440001002000802880040000A2020000800004000000",
INIT_04 => X"000DB0B1EC048005006002000028008522200008000004A0000004A002090008",
INIT_05 => X"1480000004000001000800400001210021200090904160000000000909080000",
INIT_06 => X"0008208504104200100000100000901010A1040145448000942100000A808001",
INIT_07 => X"04424205F0124005010C10002000042028092400884080000000020048480048",
INIT_08 => X"A0080004204840040000080A0A200A2A454002080000090A458294C240018200",
INIT_09 => X"0000000000000000000000000000007FE0614546024C1E10064251C088C4057A",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(1),        -- Port A data input
DOA(0)   => data_read_a_hi_256(1),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(1),        -- Port B data input
DOB(0)   => data_read_b_hi_256(1),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_2_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0C0400000682101010101000092D555550554161081447421116AAAAA820012",
INIT_01 => X"0A001DAAA04408028418019800610454A10E00C4000CA262012000C8A0780028",
INIT_02 => X"100400120DC92A5D044335282951264102C1C140091444504A900282D2604003",
INIT_03 => X"82921220A28080400A92560001002012E062020401AE088010808000E4110B00",
INIT_04 => X"100008000200100030000814442D54032820101802A0242A0104843012480048",
INIT_05 => X"14A500A04C448418400080141019210323C258959641002C01550509596D8041",
INIT_06 => X"80A4201F4350564188D54C2852CA5244D2A1011554501081B86100020C10D280",
INIT_07 => X"10405294C0910105021308848045913A20488481D851900022D022084AC9A843",
INIT_08 => X"A14B3D0D0149D2C08680480902A008A21444460200150B9A8D46B4AE500242A9",
INIT_09 => X"0000000000000000000000000000007FF22A53D68064DC5B30EAD404FCF071D0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(2),        -- Port A data input
DOA(0)   => data_read_a_hi_256(2),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(2),        -- Port B data input
DOB(0)   => data_read_b_hi_256(2),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_3_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C100300AE488011001100124C366666619989C84A945469141B33333120002",
INIT_01 => X"0010B50C846428208410028800800004210C0080004802E0558084412581D06C",
INIT_02 => X"1014001A2DC13AA94C09640319D2C44822849441090EA800CA208882C2250108",
INIT_03 => X"3183106A6998924449B054A0100C200804A02200110008904280808005100940",
INIT_04 => X"14000C000000108010002045042B32032829404041B00426108424284A08426A",
INIT_05 => X"0C244E664058850000200011140503090B80449596C8606070CC6109496EC048",
INIT_06 => X"80042815D38052550A05085101C3405452A1010500548530A143160258626300",
INIT_07 => X"024A001480100405020D008060418402A008060020529010218514184A492042",
INIT_08 => X"38D194A5014A7282838524114A19080AC5514649018C09AA954AACA250018A0F",
INIT_09 => X"0000000000000000000000000000007FE350C1460054143016A2C000887031D2",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(3),        -- Port A data input
DOA(0)   => data_read_a_hi_256(3),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(3),        -- Port B data input
DOB(0)   => data_read_b_hi_256(3),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_4_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C0CB20AC108100011110000100FC78787806181810800D18195E3C3C3C028006",
INIT_01 => X"081025AA604408128400100081842028A108042040C20260028008C0D4001E2C",
INIT_02 => X"920406000DD1A4110542042879D2002022409101095E64104810200892214103",
INIT_03 => X"87840669E7D0108253B6470800292C1018000000012E28885080601083130802",
INIT_04 => X"40000000000010802080000550370CA52102020207C8240E8380941A3A480026",
INIT_05 => X"0C2151E105000C211022200030214120038000919240406AE3C3212909388059",
INIT_06 => X"00806017E820421400016040008808008481421830255BA49001648258A18424",
INIT_07 => X"8048029480900024440914084041142A20480412804080801784700048488840",
INIT_08 => X"03DB9106014C4282078CE88002083AAE34F30E2B243C299A0D068C8640850008",
INIT_09 => X"0000000000000000000000000000007FED49202102283E622408110054C44518",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(4),        -- Port A data input
DOA(0)   => data_read_a_hi_256(4),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(4),        -- Port B data input
DOB(0)   => data_read_b_hi_256(4),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_5_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"CE88381F030781100000000100D7807F8048181E94A84D60A555C03FC0120006",
INIT_01 => X"083025836054C8D69416D281E46C6D2DA50DA4A0F217E665A82460C84080128C",
INIT_02 => X"918425105D45A411060604228642890040A491071E213031012C8000D7030306",
INIT_03 => X"6860699410016D322448A8D206009113042000042000102A0082501400108001",
INIT_04 => X"55FFF3B1EC0794AD34E02A000040FC8440091018B802AE516C689E45835CB911",
INIT_05 => X"30000C134C5C8880246048952206220929040520221628122C3FA5920220C049",
INIT_06 => X"86ADEA0D46F084351A5B0A506EB686DD148BD0C23D133042100590000000803D",
INIT_07 => X"0AEF157C82B90406B1CD3000653D617FE15C8680B883100328628A1890833CE4",
INIT_08 => X"542D8DA40091A20280520C894A111048030004C0B34352B41A0D190C8001817B",
INIT_09 => X"0000000000000000000000000000017FF07800000EF9FA8F76FC3ED7FDBCFDE9",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(5),        -- Port A data input
DOA(0)   => data_read_a_hi_256(5),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(5),        -- Port B data input
DOB(0)   => data_read_b_hi_256(5),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_6_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4CC0718E26481111111111000D7FF80000FE01E102005601155FFC000000002",
INIT_01 => X"0810258C61440802842102C018619210A10840B00C14B062001008C094001C2C",
INIT_02 => X"120420000090A4110402042000420000088091010002201000200000D0010102",
INIT_03 => X"400010080000000208505481800020D004200004000208000082000000121000",
INIT_04 => X"5400000A10C01088B08168555508028528010000000024204000842102480108",
INIT_05 => X"040008014404088003000604220103210004009594C000024000080959480049",
INIT_06 => X"0084200940205614084100400080800004010000695C48419401100000008000",
INIT_07 => X"800800148090002445090008400100022048049210518081000404004A480840",
INIT_08 => X"A0098004014852138806E8810020080201000E032400299A8D46ACA650850008",
INIT_09 => X"0000000000000000000000000000007FF83BF7F7867CEE7F72EAD507FCFC7CF8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(6),        -- Port A data input
DOA(0)   => data_read_a_hi_256(6),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(6),        -- Port B data input
DOB(0)   => data_read_b_hi_256(6),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_7_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4CC031862648000000000000000000000000000000004000100000000000006",
INIT_01 => X"080025A020440812842112C012099638A10044B009001060000008C014000C2C",
INIT_02 => X"100400020080A4110542042800C2040000809100000220100020000090010002",
INIT_03 => X"4000100800121818484010808040085024200000012C0081D080000000100000",
INIT_04 => X"00000C04120809004010C1000028022009090000000065204001852102CA0428",
INIT_05 => X"C82948000444A41041208215901060020B82100504080000400004A040570400",
INIT_06 => X"0180213F99301D00804044404008800014010800544010411001300250208000",
INIT_07 => X"1008001481941105010910044040100820CA0C81881900018004021002020A51",
INIT_08 => X"00026005010011C102040028081810841500000002000000C060202010010000",
INIT_09 => X"0000000000000000000000000000007FE2000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(0),               -- Port A write enable input
DIA(0)   => data_write_a(7),        -- Port A data input
DOA(0)   => data_read_a_hi_256(7),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(0),               -- Port B write enable input
DIB(0)   => data_write_b(7),        -- Port B data input
DOB(0)   => data_read_b_hi_256(7),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_8_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"D08800000008000000000000000000000000000000800C000100000000000002",
INIT_01 => X"081425A001440802842002C000090410A10800B000140062000001C80080000C",
INIT_02 => X"100400020010A4110542042800420000008011014002200400200000C0010142",
INIT_03 => X"500000080802020000584481840028D204200004000208008080000000301000",
INIT_04 => X"0000004200002040880B00800000020120010000400020005000800102404000",
INIT_05 => X"8400080044040000032006040003250101000191904200805000001909880010",
INIT_06 => X"808400050012420508004840000A804404000001200000409001300000008000",
INIT_07 => X"00080014808000040109100040401000204004009940880110040648C8D92800",
INIT_08 => X"4014190501CA5011880400010200180E010006400200191A0D068C8644210000",
INIT_09 => X"0000000000000000000000000000017FE74B67630200DA6122CCA8C0FCFC7D61",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(8),        -- Port A data input
DOA(0)   => data_read_a_hi_256(8),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(8),        -- Port B data input
DOB(0)   => data_read_b_hi_256(8),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_9_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100204811111111111000000000000000084084C008100000000100002",
INIT_01 => X"000025AAA0440812840112C000609228A10044B00000B060000008C014000C2C",
INIT_02 => X"B20427820090A4110542042801D2046008C00000010264104A302002D2214003",
INIT_03 => X"5000100808000A100850448800202C1014200004012E088050827814C2B20003",
INIT_04 => X"54000C0002081088308028555508020120090000400000A0500010A102014008",
INIT_05 => X"14214803445888001000201120052509090004909250088250000DA909BF8459",
INIT_06 => X"8024488D001242050A404840400A825400004411090100409401300258208000",
INIT_07 => X"020A10948002C4244109100040401108A0016610A942908020040258484B2008",
INIT_08 => X"200000270049E000800404814030080A00200A402200092A158A94CA44210003",
INIT_09 => X"0000000000000000000000000000007FE4234A4E04D5408102225FC4FD58D982",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(9),        -- Port A data input
DOA(0)   => data_read_a_hi_256(9),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(9),        -- Port B data input
DOB(0)   => data_read_b_hi_256(9),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_10_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C4C800100264811111111111000000000000000084884C008100000000100002",
INIT_01 => X"081025A360440812840112C000609228A10044B00000B060000808C014000C2C",
INIT_02 => X"100400020010A411054204280152000000801101010220104820000090210102",
INIT_03 => X"4000000800000810004800880020040014200000052C00805080000000100000",
INIT_04 => X"54000C0002081088308028555500028600090000000020004000800102400000",
INIT_05 => X"18214802045C800010202015000642080900050102980800400005B01037C449",
INIT_06 => X"80A0480500200401020008404002025500804001010000411401300A58208000",
INIT_07 => X"024A101080800404020914804040010080400600300310012004041880932800",
INIT_08 => X"400000270081B01000040400423010040100040002001030180C180C00010003",
INIT_09 => X"0000000000000000000000000000007FE771F0778E5016F81494EC15A01C5DA1",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(10),        -- Port A data input
DOA(0)   => data_read_a_hi_256(10),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(10),        -- Port B data input
DOB(0)   => data_read_b_hi_256(10),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_11_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C2880203B0600020202020200000000000400000000004001100000000000006",
INIT_01 => X"0824250C40448882840602C168004100A10180B0B4004064000000C00000000C",
INIT_02 => X"1104001010042411060204000042010000801104540220240024000080010042",
INIT_03 => X"40000888000041002040009302000181042000000000000A8080000000100000",
INIT_04 => X"006AA26948820D258C10C2800000020000010000100000C0402000C103962001",
INIT_05 => X"800008000400000006400C800000000001000000000000004400000000000000",
INIT_06 => X"0401030500000000100000400420000000029800000020401005900000008015",
INIT_07 => X"80840508832D00002489200840184014419604020000000000040000000012B0",
INIT_08 => X"4000040400000010000400080808008014000000120020000000000000850300",
INIT_09 => X"0000000000000000000000000000007FE7394D4E04C1148010440605A158D940",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(11),        -- Port A data input
DOA(0)   => data_read_a_hi_256(11),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(11),        -- Port B data input
DOB(0)   => data_read_b_hi_256(11),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_12_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C88A1F83F000020022002200020000000040004000000480012A000000000002",
INIT_01 => X"081025A00054C8C6940202C06F000801A50080B037810465AA0C60C00000008C",
INIT_02 => X"110400125014A4110746042880428100008411010603302100248000C0030106",
INIT_03 => X"4000018800010400044000DB822095C1142000002000102B8080000000100000",
INIT_04 => X"01F36369D0410025CC5281000040020000011010200000904800008103978000",
INIT_05 => X"E00808004C00000037406E800000000101000000000420004800000000000000",
INIT_06 => X"040D038504000000180002502604008800029C02000000421005B0000000801D",
INIT_07 => X"00000400832EC000820D248065300040019764000000000280048800000012B4",
INIT_08 => X"2400040700000001800400010000000000000000024000000000000000018060",
INIT_09 => X"0000000000000000000000000000007FE701B2B18095005C029A931235189910",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(12),        -- Port A data input
DOA(0)   => data_read_a_hi_256(12),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(12),        -- Port B data input
DOB(0)   => data_read_b_hi_256(12),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_13_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C6CC00100206811133331111580000000000010084084480A320000000100002",
INIT_01 => X"083425A020C40812840552811060DB28A10144A08801F060003809C014000C2C",
INIT_02 => X"114400321014A4110742042803520800408011054102201449240000D4210342",
INIT_03 => X"4800000800016D300048A0880020041014200001832C10A85080020000104400",
INIT_04 => X"559C5DAACECB908DB8EB6AD555400212408901093800EB004C298B010240A800",
INIT_05 => X"0821480244D88004304060910006428909000521229208014C0085B21237C44B",
INIT_06 => X"03ACC805002184000A1002402434028800004002008000411001B0065020801C",
INIT_07 => X"0AA5156880800412B2C9048040306145C04006083083104128040C309092080C",
INIT_08 => X"C00004270091B0008034044140101044020004801A0052341A8D194C82110153",
INIT_09 => X"0000000000000000000000000000017FF83800001EF9FE0F76FC3ED7DDE4E5F8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(13),        -- Port A data input
DOA(0)   => data_read_a_hi_256(13),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(13),        -- Port B data input
DOB(0)   => data_read_b_hi_256(13),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_14_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C088000001600222000000005A0000000040014000000480012A000000000002",
INIT_01 => X"08002500004408028400828000600000A10020A00000A060000000C00000000C",
INIT_02 => X"1084000000002411040204000042000000801100000220000028000081010002",
INIT_03 => X"4000000800000000004000800000000004200000000000000080000000108000",
INIT_04 => X"0001B0E620C72800004202800040020000010000000000004000000102000000",
INIT_05 => X"0000080004000000000000000000000000000000000000004000000000000000",
INIT_06 => X"0000000100000000000000400800000000000000000000401001100000008000",
INIT_07 => X"000000008000000000090000400C000000000400000000000004000000000000",
INIT_08 => X"2000004400000000000400000000000000000000020000000000000000010000",
INIT_09 => X"0000000000000000000000000000007FE07BF7F78E54CEFD36FAFD17FCFC7CF3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(14),        -- Port A data input
DOA(0)   => data_read_a_hi_256(14),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(14),        -- Port B data input
DOB(0)   => data_read_b_hi_256(14),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_15_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"C08800000060022222222222000000000040000000000400010A000000000002",
INIT_01 => X"08002500004408028400028000000000A10000A000000060000800C00000000C",
INIT_02 => X"1004000000002411040204000042000000A01102160220000020000080010002",
INIT_03 => X"4000298800000000244008800000000004200000000000000080000000100000",
INIT_04 => X"0000001000008564843100000040020000010000000000514000004502000011",
INIT_05 => X"0000080004000000000000000000000000000000000200004000000000000000",
INIT_06 => X"0000000100000020000200400000000000000080000020401001100000008000",
INIT_07 => X"0000000080010000000900004000001000008400000000000804000000000000",
INIT_08 => X"0000000400000000000400000000000000000000020000000000000000010000",
INIT_09 => X"0000000000000000000000000000017FE0000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(1),               -- Port A write enable input
DIA(0)   => data_write_a(15),        -- Port A data input
DOA(0)   => data_read_a_hi_256(15),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(1),               -- Port B write enable input
DIB(0)   => data_write_b(15),        -- Port B data input
DOB(0)   => data_read_b_hi_256(15),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_16_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"05104816EA00C199999999998B82D55555055577C0000675C3816AAAAAB80003",
INIT_01 => X"8014102000081213688B1862C400120ADA22C61962221218A90010E0957F0E0E",
INIT_02 => X"C200BAC50001061C8901300A2C0980A50085C801003641100400A00980206443",
INIT_03 => X"E2D5423CB284889002E20281C02900E8CC00000340A9401040162E6680824001",
INIT_04 => X"FB58CA2929ACA9E021F940410505564001B30303829FBF0A61DAFF19988017A2",
INIT_05 => X"C02C5CB08D408884438B07110220080204209000000028BA6155252000033165",
INIT_06 => X"2420A0A00A840000022800281241080040000208000005E4321254B281295280",
INIT_07 => X"2200000001020208023485003A048820088005000200124342D6311100028200",
INIT_08 => X"91612A8AB000AC00B4C661304000200000110027431500000000001000005485",
INIT_09 => X"0000000000000000000000000000017FE0334A4A0C60F6FB363875D4C538399B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(16),        -- Port A data input
DOA(0)   => data_read_a_hi_256(16),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(16),        -- Port B data input
DOB(0)   => data_read_b_hi_256(16),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_17_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4F74BF57E6E587FFFFFFFFFF92D71999998E665DC000E1D9E8758CCCCCF80000",
INIT_01 => X"2ADE30F033C915094A13393EDEF4B2265284CE4B6F40B85001AE0AB1FA003513",
INIT_02 => X"664123B786736A3991E3A47C1D59727F83855D59A1AC21CA6C30AAA2F8F149E3",
INIT_03 => X"01EF407061DE98DF4182021FC45117E22A0888D2C6F8E0FE6823B275CDE77725",
INIT_04 => X"BB2150ABD272C2B36B5D7FAEEF833D7807BE272701DDBF0600D8FF080FE617A2",
INIT_05 => X"00F1B07EFE79DF5FFF8BFF72DD78043DCFAFDA000117AD7600CF4E60001399BD",
INIT_06 => X"3AFF5F17BF430142FF1415AD12C11700001FF800FCFF5D0421B948FFE3CB1CD7",
INIT_07 => X"77105801B3FDD2780225C3B59F058DB28BFEEC394102168741D8107700029BCB",
INIT_08 => X"A0E66D1FC40024DFE9C023F3F007600088771815600D0020100800010630ECAF",
INIT_09 => X"0000000000000000000000000000017FE00C363180DDE2F82193AAC100343592",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(17),        -- Port A data input
DOA(0)   => data_read_a_hi_256(17),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(17),        -- Port B data input
DOB(0)   => data_read_b_hi_256(17),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_18_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"80900040060040000000000040039E1E1E0F80060E1C067E2F81CF0F0F000003",
INIT_01 => X"82500F0000100211A6110064200002886984501A10005048A99041D0557F0A28",
INIT_02 => X"C0404B0000108804C04211220424A28000C0804940226454001080009001A502",
INIT_03 => X"6078001C3080000000EB02801129001CDC40000100810011D008380302004002",
INIT_04 => X"14CC5F2ABCE128A014BAA8011400FE0280431018808040026081000988000002",
INIT_05 => X"CA0C5C1101DAA0A0038007000206DA400000054342A00210603F31943425E248",
INIT_06 => X"3520A8A040AC0C8020A920A081014C00C208070C000001654B10548004316700",
INIT_07 => X"00005000000104000A360D0295820000000082043609210080661584A1B44430",
INIT_08 => X"90266BAC10A190201046240000001405208005018303969048A41A4C084AD080",
INIT_09 => X"0000000000000000000000000000017FE00917109AA06CA940889D014484C5D9",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(18),        -- Port A data input
DOA(0)   => data_read_a_hi_256(18),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(18),        -- Port B data input
DOB(0)   => data_read_b_hi_256(18),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_19_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"00014020080007FFFFFFFFFF82D7E01FE008005FC000E7E1C1F5F00FF0380003",
INIT_01 => X"0000000000000004108800000000000104220004006A80000000000000000000",
INIT_02 => X"00009440000005400C0000020400000000000000002200000020000940000000",
INIT_03 => X"6040001C3080000000E20280000900000C000000000000000014440010000010",
INIT_04 => X"0031E06403EF80AC801BC19055000E0000030000808000026080000988000002",
INIT_05 => X"00001C1000000000000000000000000000000000000000106003000000060448",
INIT_06 => X"0000000000000000000000100000000000000000000001641063748000048020",
INIT_07 => X"0000000000000000000000002000000000000000000000000046100000000000",
INIT_08 => X"9021104020000000004620000000000000000001030100000000000000000000",
INIT_09 => X"0000000000000000000000000000007FE02EDADE84C87AAA0501480081CC8CB8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(19),        -- Port A data input
DOA(0)   => data_read_a_hi_256(19),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(19),        -- Port B data input
DOB(0)   => data_read_b_hi_256(19),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_20_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"00000000000007FFFFFFFFFF82D7FFE0000FF85FC000E7E1C1F5FFF000380003",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000027C00000180004400007E00000000000000000000",
INIT_03 => X"E7C6867DF780000093E60380000900000C000000000000000000000000000000",
INIT_04 => X"5402305271203D4CC80008550017FE000003000087E2008EE386009BB8190046",
INIT_05 => X"00001DF000000000000000012000008604008000000000F9E3FF000000802803",
INIT_06 => X"0000000000000000000000000000000000000000000003E40000548000000000",
INIT_07 => X"0000000004025200000000000000002008012D000000404007E6700000000000",
INIT_08 => X"33E0040100040C4805EEE00000000000000000230F3F00000000001120000000",
INIT_09 => X"0000000000000000000000000000007FE0402621121D803000120200200848E0",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(20),        -- Port A data input
DOA(0)   => data_read_a_hi_256(20),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(20),        -- Port B data input
DOB(0)   => data_read_b_hi_256(20),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_21_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4410801502168D555555555520D7FFFFFF90001F8000057F8D55FFFFFFF00002",
INIT_01 => X"8880BE000439376128C090A2E09240284A30242970600098540084F0017FA04B",
INIT_02 => X"0511481A600817F8800B64437D11428202208800047EF900C80488000085480F",
INIT_03 => X"E7D80EFFF7CC20E513E60BF2044D11000C800040108C0022022B789ECAA60068",
INIT_04 => X"54672E114C020425140002000017FE00050366668780201EE380801FFD140436",
INIT_05 => X"00801FF2120218A12488494149C000200840400200040578E3FF002000170449",
INIT_06 => X"4401A20026C000403008142D00504C00C20E9308545453F43B10568027417811",
INIT_07 => X"1021004806380400821589B43102800083140200010000811FE77000010054A2",
INIT_08 => X"DBF7F9E20001A3C285CFE02200024000A2D500B307BF0020100800000000F056",
INIT_09 => X"0000000000000000000000000000007FE038888C1EF9FE0FF6FC3CD7FDFCFD78",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(21),        -- Port A data input
DOA(0)   => data_read_a_hi_256(21),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(21),        -- Port B data input
DOB(0)   => data_read_b_hi_256(21),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_22_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"6CD0E84501520D555555555524FFFFFFFF90009F8001C17F8055FFFFFFF00000",
INIT_01 => X"0A94BEAFE77D3C314A43D337A45241685290F4CFD22090F85C488C03D57FAC62",
INIT_02 => X"F6157F9A78589FFDD14B756901537001E028C4415900AB14E83DA22A50A5694B",
INIT_03 => X"0827A802001090086000807A1124150890A222023DA002AA52AE78DFEAF6314B",
INIT_04 => X"55F76721460910AD34C028555540006045287676087620400446A00045541AC0",
INIT_05 => X"00A54202485AADB1748AE9510DC4080B28684420220661000000F582022384C9",
INIT_06 => X"54ADCA00000680303A0700FD92A012001036D0C05454D0103B30222A055BFFD5",
INIT_07 => X"1284170066A90561124C8480FA0545630B5480B00288111730018150100258E0",
INIT_08 => X"A817FD23001023D3900105A3409342604044500400800084422111088C6164DF",
INIT_09 => X"0000000000000000000000000000007FE07B77739EF5EEFB76BAFF15E4BCFDF3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(22),        -- Port A data input
DOA(0)   => data_read_a_hi_256(22),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(22),        -- Port B data input
DOB(0)   => data_read_b_hi_256(22),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_23_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"8A99D0720284A800000000006A000000005FFF400C1804002D00000000000002",
INIT_01 => X"A00080000420E3E7BC8241B640909201EF20906F206006E5F4E2B4F0200040CD",
INIT_02 => X"A39050087D451C8190084003FC04B16802C11910167EDC8180382AA20006800C",
INIT_03 => X"E7C02FFFF780000017EE0BA0044D00122CC888D0700CC010020D0094F2A38B73",
INIT_04 => X"019955B0C4038005006002000017FE020003404087818A5FE3980A5FF8000017",
INIT_05 => X"08001FF91300365040888000D01242000282110100900878E3FFF03010124000",
INIT_06 => X"320820000420040000B034B10850100000010004000027F510105680275BFFE8",
INIT_07 => X"000000000000100002134014B008841000000801100108000FF7F40080908000",
INIT_08 => X"1BE000800080100005CFE00000001004A091043B97FF1200000008000002F834",
INIT_09 => X"0000000000000000000000000000007FE0000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(2),               -- Port A write enable input
DIA(0)   => data_write_a(23),        -- Port A data input
DOA(0)   => data_read_a_hi_256(23),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(2),               -- Port B write enable input
DIB(0)   => data_write_b(23),        -- Port B data input
DOB(0)   => data_read_b_hi_256(23),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_24_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010800820001080000840037C00000000000000007E88008380000000040008",
INIT_03 => X"E7C0067FF780000013E603A0000D00000C800000100000000210008001000040",
INIT_04 => X"000CBCB020070000004002000017FE00000340408780000EE380001BF8000006",
INIT_05 => X"00001FF00000000000000000000000000000000000000078E3FFF00000060000",
INIT_06 => X"0000000000000000000000000000000000000000000003F4004C568050200000",
INIT_07 => X"00000000000000000000000004800000000000000000000007E7700000000000",
INIT_08 => X"3BE000400000000005CFE000000000002091002307BF00000000000000000000",
INIT_09 => X"0000000000000000000000000000007FE01D1A18B4B598CC60523ACB39BEBD60",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(24),        -- Port A data input
DOA(0)   => data_read_a_hi_256(24),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(24),        -- Port B data input
DOB(0)   => data_read_b_hi_256(24),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_25_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000D555555555524FFFFFFFF90009F8001C57F8155FFFFFFF00002",
INIT_01 => X"0000800004202020000000000000000000000000000000805400840000000040",
INIT_02 => X"0010000820001080000840037C00028600040000007E88008000000000040008",
INIT_03 => X"E7D8067FF7DC38FD53E623A0000D00000C800000100000000200008000000040",
INIT_04 => X"00000C018C008424042000000017FE00000340408780040EE380041BF8080426",
INIT_05 => X"00001FF000000000000000032224042808040002000004FAE3FFF12020B68010",
INIT_06 => X"00000032FBC009428008000005014C00C2080308000003F40000568000000000",
INIT_07 => X"00A5414910100400B0C0092001022015C00802002102008007E7700001000403",
INIT_08 => X"DBE002201C05A0000DCFE00000002000229108A327BF0230180C100C00000022",
INIT_09 => X"000000000000000000000000000000FFE020272920E9ED0B200C52CF20B83A81",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(25),        -- Port A data input
DOA(0)   => data_read_a_hi_256(25),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(25),        -- Port B data input
DOB(0)   => data_read_b_hi_256(25),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_26_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"85F820440E61E5DDDDDDDDDD81D7FFFFFF8FFE3FDEBCEF7FDFD5FFFFFFF80007",
INIT_01 => X"AA5E3FF033CC1A1BA4993AAC8064328EE9265EAA400ABA7000401AC1DE00573E",
INIT_02 => X"F645FFF78F73EF7DDDE3B57E7C6F72BF89C15D49E0FE675E24302AA9F8D1E5E3",
INIT_03 => X"E7FFD67DF7DE1ADFDBEF578C5479263E7E600053CEFDE25C78BFFE7FDFF77F3F",
INIT_04 => X"FE000C000338529A33843C7FFFBFFF7BAFFF272787FF302EE3D6F03BBE6057EE",
INIT_05 => X"0ED5FDFFF7FBFFFFD889B133FFFFFFFFCFAFDFD7D7FBCFFFE3FF7FFD7DFFFFFF",
INIT_06 => X"38F65C3FFBFF5FD6EFED75ED91C9CF11D688635CE8EB4FE5FBFB7CFDF7FFFFE6",
INIT_07 => X"77525A85B4C017794B3BCFB7DA839D8AAA600FBDFF5BFFC567FE77F7EBFECD03",
INIT_08 => X"B3FFFFFFFDEFFFFFFFEEEFF3F2377C0F29F31F676F3F9DBA9D6EAEBF7E7B7C8F",
INIT_09 => X"000000000000000000000000000000FFE0034B422CD53444E373420BBD2C2CFA",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(26),        -- Port A data input
DOA(0)   => data_read_a_hi_256(26),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(26),        -- Port B data input
DOB(0)   => data_read_b_hi_256(26),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_27_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"11200008002844CCCCCCCCCC80D7FFFFFF8FFE1F5AB4AB7F5ED5FFFFFFEA8015",
INIT_01 => X"080A0E5012800008002029000029049200080A4000142822000002090A800110",
INIT_02 => X"4441D8370DC3416110A004547C8854AB88011100A0FC000A040022202A1000A0",
INIT_03 => X"97EF9671EFDC1ADDDB97570404512A062A000057CA7F0844783D024B19456E38",
INIT_04 => X"FE000C000338529A33843C7FFFBFFDDDAC8E252547F7102E93D6603A3C2056EE",
INIT_05 => X"1611F1FEB2FFF65648209017D9D5B9CECEAA96D6D7798F7D93FF77ED6D7FBFEF",
INIT_06 => X"B0721C3AFBDD5BD7A76D7C05C1CACF55C688231D81804784CF0848A55D7E7BC2",
INIT_07 => X"D35A189424401654452153BC0AC3998AA2200B2BAE5AF54467F873BA6B6FE503",
INIT_08 => X"83FFFF31FD6BEFE677E8EF78FA3E4C8B1D1113474C3F2DAA956AA6BB7AD42E0F",
INIT_09 => X"0000000000000000000000000000007FE03F1110E441278421012A0970222288",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(27),        -- Port A data input
DOA(0)   => data_read_a_hi_256(27),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(27),        -- Port B data input
DOB(0)   => data_read_b_hi_256(27),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_28_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"4128400000606088888888888000000000000000420526004380000000080003",
INIT_01 => X"220A20501184080808802A90006000C202200AA40000A820004A02822A004110",
INIT_02 => X"B24427A5000A440440A21114001A00002288C440A980220A0CA1088828B120A2",
INIT_03 => X"0000000000008000800100041110020C8222220186D182D428827A14E2B25403",
INIT_04 => X"AA000000013042120304142AAA80013881A40303000014000000440000280000",
INIT_05 => X"02B4A005A1A149A7080A1040262094E4E444C2404123C2870000024404803B36",
INIT_06 => X"00523400000B0080050000400000110010352040D4D490005020080D02048002",
INIT_07 => X"41104A01405003310028020040000CA00828019805006CC0500800E220240140",
INIT_08 => X"400000D0E0240C34682002D2B0852621C8444918E80004004000121126310000",
INIT_09 => X"0000000000000000000000000000007FE02064636888C821822C1405C480005B",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(28),        -- Port A data input
DOA(0)   => data_read_a_hi_256(28),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(28),        -- Port B data input
DOB(0)   => data_read_b_hi_256(28),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_29_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"A5F0A0540E75C5DDDDDDDDDD81000000000FFE20C60C677EC3D5FFFFFFD80003",
INIT_01 => X"805E1FFFF1C81619E659392E8076B2AE79965E4B402AB858000A0A71FF7FBF3B",
INIT_02 => X"E240FFF78F72EB588DE1A03E016D627D81408809E0FE455E66100001F850C5E1",
INIT_03 => X"E037C67C104E00C793E9038C403806345E4000438F5D604C281FFE7FDFA35F3F",
INIT_04 => X"FE000000013042120304142AAA97FF7A87D72323807E340EE046F41B866813C6",
INIT_05 => X"0A50BC0FF5FBDBBE988131236EBAD6DDC7A78B4141B383FFE0007E541497FF7F",
INIT_06 => X"78D67417992B0592EDA015AC9001010000116000A8AB4BE16BD37C7FF5C57C26",
INIT_07 => X"75100800B0D002380A338E97988008800068051D550176C167FE04F7A0B64941",
INIT_08 => X"9017FFDFE8A4BFFFEDEE03D1B0173405A8A20D37EF00941008040A15263A7481",
INIT_09 => X"0000000000000000000000000000007FE0F480845EF1DE1EFDF8B9DEFDFCFDF8",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(29),        -- Port A data input
DOA(0)   => data_read_a_hi_256(29),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(29),        -- Port B data input
DOB(0)   => data_read_b_hi_256(29),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_30_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"0000000000000222222222225A00000000000140000000800020000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"E000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000007FE03B7F7BFCFDFCEFE37F7E0FFDBCBDF3",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(30),        -- Port A data input
DOA(0)   => data_read_a_hi_256(30),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(30),        -- Port B data input
DOB(0)   => data_read_b_hi_256(30),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


ram_bit_31_1 : RAMB16_S1_S1
generic map (
INIT_00 => X"60008010001404444444444400D7FFFFFF8FFE1F0810817F0C55FFFFFFE00000",
INIT_01 => X"08800E0FC20105004A40000200128020129000010020000800000030017FA801",
INIT_02 => X"4401D8120D410161100004407D1050EB80011110017C00804A00222200200800",
INIT_03 => X"87EF8671E7DC18DD5386030004410002280888D2492C0080503D004B19452A38",
INIT_04 => X"54000C0002081088308028555517FC40040A242407F7000E83D6201A3C0016E6",
INIT_05 => X"002151FA125AB65040008013D9D4080A0A8A140202100D7883FF75A0203784C9",
INIT_06 => X"60200832FBC40952822D340581C04E00C20C030C000007840B0840A2557A7BC0",
INIT_07 => X"1200100004001440000141B40A83810282000A21220A110427E071100102C403",
INIT_08 => X"03F7FF211C01A3C215C8E5204012400000111007043F00A05028100808402C0F",
INIT_09 => X"0000000000000000000000000000007FE0000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
CLKA     => clk, 					-- Port A clock input
ADDRA    => address_a(15 downto 2), -- Port A address input
ENA      => enable_a_hi_256,               -- Port A enable input
WEA      => wbe_a_hi_256(3),               -- Port A write enable input
DIA(0)   => data_write_a(31),        -- Port A data input
DOA(0)   => data_read_a_hi_256(31),         -- Port A data output
SSRA     => '0',                    -- Port A reset input
CLKB     => clk,                    -- Port B clock input
ADDRB    => address_b(15 downto 2), -- Port B address input
ENB      => enable_b_hi_256,               -- Port B enable input
WEB      => wbe_b_hi_256(3),               -- Port B write enable input
DIB(0)   => data_write_b(31),        -- Port B data input
DOB(0)   => data_read_b_hi_256(31),         -- Port B data output
SSRB     => '0'                     -- Port B reset input
);


end;